��/  ��^k*��A��D@7�քW�g̝�G�^�T�|�IVϪ�y�p;�5��p:#�oj#�_����슧�;|���k��I���4#�g힆D���+ؤ
OK02����l\��j��կ��wI�2W_��Ha������yf���&߽\O|Ć�Y�U����~��,��Xy7)�!fR	�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P�ﳙ�Y�+���]��%���K �ܕ'J��A�$g�k}Ӄ�l펀(�P��w�;d�L���6#S��� ( z�Pi�dc�S�t=���cWL\6�c��ܒ�uD6�/뀽��c�.���#���|����g��'�8�ڥ%�]l�Ԓ�OC#�{�b�W��>f^�Q$H�tg�{_�*���0�Io�%@��������aL�(�dU�gӽFc�_�_K�[O�✯_RpF�c��
�6˾��	�ap
_�Ժg�{9B>d�[O��H���4�ꦴ&�� ]���禺T���o�|��,�����/��5�
~���&EQ����"d�d�<�]q���]j�;�t���� ��X�Uږ`�94N!�����	Y�ˌ�\fvv���E�X�e�+0�f�,ŋ*?��v��.����EWW�dC��N��Xp\!����6���ʳV|�BR��C�=����&
7ZH�B8���K����U\��J��q�װ��'V�<��1:�'�8�G`"���k~՜_���	j���;���~}ߌ�2�Y�N��{�k&��I�Y�&�]'���5+F��e
6~��������a�
���߃	�/q�>���K𿽐`�Cm����T\��0SRg9������T�j�gܑʫ^���H����0|ց�#?�dV7x�{P^׀��$��>�}��Y+7�����#\y������Gèn ��U�U�=�����	�PKhn�e�iY��藬��d5����&&�K�Te��vB�<��F�ܲ�w�?������@����1}J��ÿR$�t��sU�,�b�.�[Xޚ����ր�O/m�� �)�XT?A,�>�ԭV�#�-W�!��Ҝ̿%A��7;����Nި����I���7s��IJ�	Tl���(�c%JZ�c�vh-��TH��%��ñ�!�M���+����7��dw����aR�H�a�f�/c3Gu1��ϰ�ⷺ��,�G��۸*�!�k��l��$��ce��k��w��?�R���F��iX�}�"��W�Ƽ�Z �-w��҃u�3�ޡ-Ci�"���"��e,�n��rvZ�2�<*D ��}���<�F���$j�W�	j1>ܴ��|*TYC�k���7��EQnt{cƭ�d�Ƈw��c=0�	7�F�ҙ�f�_0�|�>J�i���Q������&���A� �*���r��e��"���1Ш��[�)>2�3��]e(S(�9g�t�tZ6�qב6��oFΝݶ.�?�:���;ҧ���d��ٽ�S�ަ��1A0�����Z���|���6#�0�	 ��pH�=5���������L|Cude�s�z�/Y`5� B������g�?J<��4�M�8�A[�6#�EGPM�#��Tt_m�In�e9AmxT�道�O����J$�8Am��g�q������b�q��R�z�C4#�'���f�� |m�����ߓs}u��!��ƴ�BR=<pc =�\&uɒ�϶��?�:��]�Ͳ��\>����y	�}q�����g���/Ú1#n�vEt{-%Lm�D|CcQ��ź5�f�l-�������:t0u�x�o��E]�/�v6Y�c����z�8�����*}V߭�����q��]���B��v�[�̾>�3���~Yh~po�~�,�S�0��E�t�F_q�L���^V�H�")�IDn[.!�a���W��t�Y!tGMo�A1���{�䠾�枉x�T����mq�,D�����?B��K�k�ː�L��Ĺ�z�(��I���аҠZ�ۯ{c��8l��E�\��w��<D��f_��w����B�bf�b#��F�R1�WmD�|��=������!�1ܦ9���#��;�u���̕
ԩR�iI��
���4��@���I��#�k-�[5s&��Rw���ʖ�&��]	��=w
��D+%FO���N��W̨�Vf���Ie��їo���n�Ht�h �d�c��;�_�nY��&�{5�j#~�N�������c'����*��F���D&�.Y�1�C�&�f�yy%��>�K$%Q4�����f�ӊ�M�
���M.jH+�L"F�,J�L�@'}_
���6�ƣMU�ƙq��<�jrgGh@o�������U4�E��Ო���eV�VF�L�|��`�8XG�;& ��#[};4�B�{�B�
ȡ'��V�&�^J�C��)���K(�D��:��������P�I�֪'�]ֿ���W�MR$��k�V�h�L� ���֫ꜣ 8췇��{�*�C�0[>"p9$�;<�-&���>�-Ҽ�r38�o��?�<���k�t6�LU�U�����՚��C���$��\Ԡ��j>\�9�]Ov�����oOt��1e���]F�����l6��[F�6Ȓ4%�4��U����,�e���U��۝�Ţ��w����@2>0������ xf������sr%�pX��3+r�[Kn&Hx������h��.�������ZAw�Ů�.���iTMO
r�� r̆S�2K"�A�+�K����|8ju\�ϐ�ʡ� of�wM�c��ֈ����G|.�Z�@�󙴈.���Y���$U�_�us������R���p��>������,����m,��^�9H���Z�x�h��l�M��\7Bv�X� ԕ�	��O�<�q�c$�PQ�R@Z��dKm��e�H'�C`��*l�*���S)��<�0���N�'J�����y��(��M�{�2��uΧk��Rv\3��E��DO�Z.1���: 0v����>dF�������ֲ`#co���T�yz�-���5��>�=��dPp�wL�B���ST�z&w�
o7T����q*�_�|X3��>�!�R�������T�?���<�b��z�h���C�`�*T�P���+.\��Sg̲EHd3�}f�Dᎃy�W~O-����+��:��b]Ix���*3�V� �_�Ն�NL��Х T���'�b@X�Q��p=�_u.'����M'�{vӓ��_ �\��$�(�	��ޱ�)�����k� ��� q���\�$��E����'�4��b�f5����0�R5Dw�����˭���Vd�7N�"f�V�&�P�?�"�:��&1�I%
��\=���驸��3Ύ��\"\/  ��'w|�g�/���bmǬCK����DL�-�4.@sQR)N�b[m�HҧW��U�d�`��̡E�$Bֳ��YF�h7�Ӝ��o}�Y �� ߢ.�n�w��l]Tz������z
C�t'~����=5�-T���zҳ�J�Jj���d�����|~߈��xB���'���uA��U�=\g��h���'Ό�N\DDH���{�F�m��UЄ����q-��`�B>5`-,5�G*�O���oe/�jd�|�e�Z�����E�I���lh�<@H]C�-�����	A����[�n�Ҡ�����uwT����-�ťC[���ij���7E' |�׀K��t�x1�l�l(����ޅ� \y�V�"zn!j�"��	��׫?R���T��g�Zߕ�>�
�o�/k��Qrpy�$!�!� �pa�}D���%ͫ�Ӭ!|�tv8���2kt5��S�~��xsEa	�@�-M��s��6����W�����*�P�q�6f
�p��6������C�K�ork{��V|!�w��oO��W1?>� ,�,�[��~D\q�470L�iR��U��+O�K����c\<����	�Sٸ;|H{�$�h9w%���t�m[H���ρml#�bn��)���b���1,�T;����v�?��Z�˞��:�����<����:%��?(0��d)"_�S��>V�
:�`�bk�mo&��)1�*~���UM�704r�ܔ�d��3�������/.7�B��:�!���8��x+�t�J�/B�  U+&��9�͕T�]��}0S�X�W	�������Ba͏�����/A[�r^����	�	��g�_L> T	oD�*H�z��Q�N�ҥA���}��a����x��Bӻ�ݶ�g�5�� j��L�aҤ�w�H��J�v�PK@�������+�:z<��ѡ�l���2pc�`Q�*F���v�aF�L���=�*���sI�!Qb�J쯨e�Wލ;(R("�[��I>t�E0=��0��ӎ�*	�*DK�c��c�./˩e�.���`nN!�A!�&�2H���� �Щ fA��9��4f�&ʺ���
��6c�R9�ΠRymf� 8'�c���S��v"̢�3P���$�����]Ʀ�ȍ�"Nm��q�7�}��P�/%�섾�}��Du0������򏮧�O�R B6�<-�n�)��x�dwG��WMbT��X�}q�����1�X̺���-tMo��#T��c��l9�`��(iY��J�EȲ���B�b�u��-d��1�P�֧R(m���{���X�m�'����0�c^Ȉ�3��5G�b��?;%x��q�Z�����U�̔ҝF6�7y������d���՟ޜ���c��ꈿc��a��a����l�i�|և��jЊ@%Fc#iD�pZ]���L�!6,�y���o����[���G�-���[�����;ֵ	�5p��;6<Ml3��x.�f�E�c�Ԭ���h��k6��%�!�J�XҮ�%9�&?�S]�	%沦�(�M���#a���K׵-���1�b _�A6�,a�վ']��	d�_]�/LHa$$��WA��<����7;1�|h��آ
���J^��}�۞�/��H�C��Y�Ox9\��\0��ۺ]h'���r9Ie�D�����w�����xm`E�|C����������(KP�꟡?ڹ%�})��C@w�7�J�"���ƃ}�'5 �~*�R:��o�E!_��:j�c�D�@���0�k7�21�A�mm����/x\[�[�<5��DM��e�=(����#������
��3�i�����i�*����k�=���I��^}Vb4�UՊљ�^�:���ey������"P�L3{��n���[s��%��Շ���c �ʂ��Al|��@w����8���$��m��a�;�*Е�6�N�Y���$[�ڵ�*}��F��IK��k���ڊ:H�X�Κk#�.�2.��#^�-v�"�t��6C)Œ���N���Jw��%�Cmo�^{\'|5�V�ִ"i���N�������a�s���0~� ����y�~�9�
�G=���q>�|$�a�*6RaJ�P6���Ӭľv��јO��]�;���O�����<��B`
�>GݏT�A�`��B@n�6�>��v^��9��r0C(�H2����,إ_�Q\�)��QY�ϛ�x%+$	����7Vŝ�l��S�G����GU�G�^�r�׳��Ϙ�" ����D��:.��Yo�*�u��l����G���Ɓ��ȅyq�R�����d�MܝY^MwQ��9h9�vG��;��q��:���:;�u�������!5l!�1���`�'r�d|*��u����J�K�u���������ě��Vi ,Lߧ�H����Jhϵ:�[�.ۘ��� =gN�,pI�����!�1�j��	Z2|`���G�k�
!R,��`��˥�п�5qK��ެ19�Mk�^=�U�n>�w3P�z[EG�!\e3oC����m��:���~�W�88���,+M �w�o�J�P@���Ƽ���t�b��'��gȸO|ǌ���4m~��T�Ѥ'��2���9�Zr�\D�#��5ܒ�'��#f쇪(L^��#�2��+���?[ϩP^�t�5%b��.���w�8�qtjΨ�Q�Z�)\8Fm�ڻ㔨������N��xZ���Wڻ�sHA�?GK!�G�Z�5	��}�6��\.�N���x���:�@����C��*�|���D��a�H�
���M}y�\o�R���|@�a:7g�����r 쾬�-��L�O�(UC����+н��Z��n�V���|��<���&E�����Q�r&�K�rU�:�a�D��*�d)�P��Y{�q���UN7�t���ԣć�� ���S6A��ܭ�@���U-f�{oӡ<f�c�,�v���
 ��zJ���s�Y�_�F�TaĘ�l$(��
�5\�N��]h�����'��Z��2V��dD1\Ղaq�K�ω��cy[Vj[�'�7X�'��I��k��_@a���[L|H�ɠk��ٴ5�~�~�?�*"g�y���W�/=���%�~s�C��,�ٚ���E�I9<<D�z�S~��A�QE�1��B� ݣ�Ym�.�3����)��g�փM9��e�̗�9���zϪ�����aI1=�8~� b���}R���2Ͷ�aCp�?\EX��"_�FU���6C�}	JT�ܺ�Ue�_����jA}|VW���'���@��o'&=�񼹃���Vmw���x��Z���N�g�?"^`F������戮,3+ ;�b���b��%Ҍ��=���v��+�K~7Q��|=h8�i�t]�Zllѣu�{�6��>qUP�l���� �V�����N���cnxN���$b�d�!��ő���8�pca�p����Dmk�&���ۃz�J���U~A��İ`yh^���,���b����{�T�O�����\��lJW��Js%��-�p�j^�y�����7|]�q�#��s�����2� �qC�f��A�]\�-4�@�J�x���j{K���AĨ�1sS�Q5g��ѦϢ�{���ǋN��P:����-��z������]ވ!���{�Ԇ��XC:�M��_~( �,�i�SS��:���H�m�wfd��ڿ�[H|�i�P_�u����	*�;b%�	h#�Se"��C�Zˋ�B8
�ؙ��żF�*��OX�b�
�!bo��Cd.ɓܦ�����i���o"֕�c���ۉ���o���D����f�\�_�@�����8�e���ݝ�hѺ����2s�o�����  ,n��JTZY��M��\��\3����pz*����� ����Y���PYD�r$Ў��r�|h������1H.�˰�2��R�)��Ѹ�ȉ5JUv9��l7W�#�q��K�X�O@��;^��O�Y����j��v`�}��bOT��;Q�s��)�g��a�M��;!q�u���K�����#J���\vn~�~JM��q5�|��<kڨ�J���̓��k�v"��-I3_�C�Ik�����z��4J���]]�acN(��r)ʉ�Ƭ�k�2aZrmx�) ��6��[
��Q?�%1�UeC��q�>���V��+2l'r��#K9���se�?0�[�vi�hO�9�ҼIz�
�Cw�o]V�`賽��:��A���D7�T~S&���8��<Q'�:��0|7g��)=pƀ��7K_��`wD���lA3�l�+���5,B�mF��o����B�8g�����\���/K��P6Q~mk�Koe�'Pv�!��,	K3��M% �s?�5��s�[�U�\i�\�-��[�$�b���&��K�dT�ꑄ��)R�:�')G)x9		sc�K��m�������
���">;b���yw�#=��9�s֤ǳY�Bk��'��3̴水LR2�:jS��ޒ��-�	�<��Ǭ��f�ҏ~�8���S�L��m�v�������ze����`�⹚)@��W�5�cxg4�g �WHAo�!6�������x�L�pXh�]����b)FЮ�s#���9:�~�g�	���r��A%��̑�d
���-۴Q�-)ù�O�x2���d�Nr���)����nN��W���b�V�TKoԌ����� y����.SH���}�~]'�YL����{�kL8��y_�±���|=��Aۥ��x"`h%裞�Ź[����B�a�����[��;�� yĝ�X��\T&ˑ{�����9ii�á�y�+��0�V�C��	&<�� 8H:��8�2^�i0dG_(`(� b!e�8��Y6�p�٦"���},u�$�����KF�:4	�X�w�p����3��< �ζ��o��-7Y� *g�*DM+�a�V�:����Ma�HY�ڵ�=������g���M^>Q]L��<F$H?pP�bW�g���8u��h2Ap)�1�c!A�5]������fX�{�S�fצm*&�+[��+D>��b��-	^�{�ꖶ���f�I�ķ��3*%X{�K��:����
(�CǓ���c`�+�"c��Ԗh��U
������?[�!���`I>�Ϝ��}�	��f��`p���pl���֝�g�r����pi�^G�8�ۅ��q�rQ"�_��x���j��`�2�*
Y��T�ʭ1ڽP�'��%&k���i��
��oOy)���M�RJf 9�]��E�Ã�R�T��P-e "���j�\\}��O2,j19�#�Fj/��G� \9U��L��Z�#~��v��,tL#��ά�\��?IqZ���|J�CZ���3�#�\��pM@{86�9<r}ӲYI[�t?!#؁A�I��Q�#P,��$��l ow�`MV��~$~B�_S4�J���@��"y���XC� 
� ��+9IG_���.�t�A�R��R"�v�Ah���I�H&�2]Ը�ƾ���p7�e�^�L�5����$	�+�1ނ�A������qm��h�l3�vܪ	c�h����<n� @B8�Uu����֒#XH>t��z�0a~��0t��z�VR�3)���슑�7���>���y�V��u��3{�J�G�Dy�8:��N��޻XLhEZ�f&'T$�/�vj�=�n���D��DpB@q\%Et�'�_�+�;�<�W������E�xt
;p���~�/�%y�w�qHb�d�d���1B�l�ż�.� L�"�R���c�!����Ӯp��IE���(  %��e���T�k[��5�~���C����ቸ$(��K�T�+Ћ]�����q��m�M���f�HD�M{����Rg㿨���_lo ���DH~=�_��W:+��1�P�"����jbx�X��r�ĵ�ǵJ�O�j3.����`t���{����K���۷b�- ӊM5ɇ��� �@���C@-�����nC�pԐ	1m�\�˶�Z?��h�rk��}M�v�=��h��=�X��P��[6~�6�0��#텽���k����i8AKN�:R�qqGʈ�!�ۃ�4��CEM�Y�(��0uD�Lf�����$&9f�gЁ0k��G�&�i�~�kL�0P-��@�z,�Ӎ@��*z I�L��������N�-�݅;�����H�B��� �#���+�ɲ3�Y�{x�����e�Y�uD�=q�W$s'ˢ��j_ǆ$j�c����g�OZC�ʢ�˶~����# �A��QS�w��vZ�pv�UÆ-X��&8�ҽ^cKB�W�UX�+��b=�w�����W4<8фI�~�n�<�|6��X_�g�����k�.��8_����#u#���	@�Jh.��{��2A�W+�tT��T����V�*o�0��6�&�f����'r�H�`^�;頻��Տ"����5 ��A�Mt�u!zz��>x��{n�z􄾧�݋ o���i�PY�L}����ޫ�a��$�k�8f;'�FG���P���)��)��?fI���(om*��b�7�>�|�711\6��|��� �.�u9�x�}�kR�D�5`��PsC�^�MP�i�M#)ѱ:��na�u],�2�M*݇oz\�AVv� �E�q��
%�P?O<��욂X4> h���0f_ܿ�҆�:^�2�
`x��Љ?!�%t���m����Qꋼ�$M5f�%1��n�.E��4A�ܼ�k��7�nM�_0Za�CO�i끿r����Qt�ݑ;qn?�1έOf�U��Q��<�ќ2�~�؏gR1j����=�I8���0t����CŸ"F���>���.GI�'��f���w$Z�Q�dyZ��U�v/DX�U�i�';\���5��ٍ�쭒7C�J�V~��
u�Φ��Q�e�Td���y,H���*噸t%��쫏j-F֎�SS�Ԟ�=����{f;��~�l���G�:B�wa/�+�t] W�V+��l6�Z&��fʡ%�z�_(�����63�����I�1ߤ�wa�)fGo�5C�y�HM��lCKm_|B^i+��F����ul8ލЮ3�#��w�}��1�#��rܬ�������@�l0��"���ũC�����!B:�P��$"2M�;�dI�|l�xdgE��[A�-��>r��:3�Qk�7_�`e�������S�͠�\�_�����;o_��M����0V�C.�M��@���G�R��?�j�I����F�:�M���u���9�S����l�cW,G$wDګT�I�·�	��p��Ԛ�*V\�Á�5gxǦ�i�H:�mv�o�����Oc8�jbż�]�@c��2�#��b��k?�[v��c�����o��+z�c�������zi�3)����%)�Fr�t�׿�){����3�+�JNTs�:�'0�'5Ў���u�lG��a'��r�!Z�Uz�fV�;�|9�[~�p'��A�����p�"}"�H��Sۙ6�v��TbKͿپ�JP���EV�]��P�6x�����dn��V�����I�u����rZ�(9�+��>6D� -�� ��<�yEqpZ�\�A�]�	`ޅ'Ґ�V׏������XC�fu_����L:�����#BR�P5\m)��?c�<*��W���f���)�r�x���'TE�w�.]����M�-7�W��7$��H�C躸7�u�u�4Q	VzA�>�b3�9ǃ��5;�`���MW'Wʵ�����NulQ�ݮ���u���M`Ɵ\ή�:Ux�ێ���	�t���}&]}o �!�#�c"pݩ5�}/�e'� (��
!�ؕ1�����ZDt�pL�h:@R��J�̰D�YX�He�N���5VYL�g�5��c�oc+U
Q��kg8�����]����"�@�D�ۢ2�}LŖ�rY	�����ܮ��($B�G�;ۇ�}�  �5D�����<2��oM0*� uL������w�GpL���PFvC1웰Ws�:�J�M���UA?��l若�Zv*{;��I��v2̳4v��Y����r'rnv�LXY���Ur���e�p�
����n�bVD
:�+W���g"\�S1�"���;���I�	��⚂�v�Ӓ�t����`�k�qa4H0�ꉂ��j��!�ߘ�
G�C��ѤF��oQ�W�\���:j:�k�sw�)v�� (q��X�sOO�zr���YеK�X���u��i+=��+2��$�0��}��E&=���ވZs�E)/B�\�Tv�2=v��O�G'�Dx�h�t�IUB�rh� ӫ���/��'OL���L�;�P%�T�S�.����`��59Xj�O3����~��#˝���%��G�K�r�=p{/�zw���B-�4fh=^�~���*?���l
`E�
�`����ҋ�����b��	֢�߭�=r�x�N��Gŵۣ��?�d+@s#��
�Õ���F��@!�����	�˶t���%v��M�֎���y	���ހT�創�׿�(c���9��B�S�]O)�k}$���/��8���#��"i<f]��7v^Q�R�|��=r���q���H�|�	^�.���~�L2�P:�fӅ��� ���_�l	�i�����,/�710��b(wq|d���@-f���N.�X�P��rw5�%�����E�>+�$�f���E����$�ǳ����W��LHi�J��y��eY��W�[������z+3gф�b�=3Ά��W�a>8�C}����V�)&�	?� VS�KSh�Z3z5I���n�*�%[ꄂzEY����P����Ր��k0H
�~+�JI�h�"��ƛ�����zp��2J��6�'J�u�A �*�۾��2���%qfj�1�u��XE3�����&2�2�m�ы��ʴ:�B���H�tɰ;�]�����Z@/�G�'G��1��5���#�O>y4��N�/W���xQ�Wܜm#��@j�5��,�Qݛr@��q�΋�SF��ڳ���o�qVPñU�¿�++���|��f1)�yZF��G�Ђ��4��}o���:����$�;��ǗL[eʩx�f{4b��B� X�Ir����箚��I�E._|��+{�^��� ���_M����pr8q�ȑ����Խn�2��[}t�x��tm�E���r_߇�o�lK-�%�	p�,���ֽ۷�L+ew�o��XР$XbR��ꌽ���{X�;�-��w�v�qƮd��J�֡�{V!��U�=��v۠��}2~���^㾪��t��6�R[v�k�ˈ��t�k�\���1Lt���҈qp41���o���\5����R:$OӚ�LZ�5��Ny��Z� 汏Z^���i��:c6���|;���%[�c��v�����'�	z��T��Mnֽ�
���V��9�x��R	�ߝ-��}q?�oک��ϸe�l�ל1�:-ɐ�i���h�1��+
�	` �k����T����Яf�.�!g#iA;��i]ާ8>?8'�t��KZ�����N����>�_Y,�(sy���Ῐ�Fn*�xA�ݠ���Zњ������j�yA�f�Ȧr�5���.s�����9�Y�^S��H�����M��%���H�e�ć7�GІ��rc�#΄�ć5�|)K�F�zj�`EKs�w��X����ˢ��%S=����.-"n����K.�U*>m�+o+�ɶ�yme��(��SZ�G�_�R��9Э������$�i�pX�~?�;�4�q�śwG����&��+���$�/�Zx�)ߨ�t]ς+op���<dX��t�&��șQ"��E`87�dp��:7l^&����>J@�	��N	#Y�ݓ�_<�Ap IgB�+�r�d^���g�2>��a�W�=M��W(����=a���@Fr��G\:��@D��_Hd�ֆR'k7eH�)��E>���l��E)�wD�겼'��_��3Qj��+7/M���T�j:���]�6Q���� ��&�d� S�&s(Ģ�C`��F�ix4�,��b) �V�nU~F�s�u��zP�y��ʡ��d�0]�?���'������n�xt붡��쫙U�"�1 ^bF.�P�!��0B�UC���j�^:n�'cZ����w�P���;�7��NC��)��V�ѽ�H��Q�Y�b �JVL�"�����l�x2Z�MV����d`�Z�Ckα����Ԡ/��3�ިL�r�^>/i�B'��I6>��zW#2���(�,����\hl���J!�Փ��ŗ��uV�G��#�Nʤ�����0VzH%�K"u����5Hp�q�85�놐V��Px$�4���ʽ����X��c��}��n=ݳ=PuG,�9� �A��@G>y5L���Ҳ����4�'y�.Lr<U@k��W�]�C�M��2k�fn�hj4}��L�[#�i�"��s����4���������B�:8���b�f��%.�%�Th:��i���-�3%��1�#<��ts����,�3�2��[}�TkՖܕ�S� �'�K�	:x���sg����d�ƿkio�~
_�]'z��
�/4�����R��}9�Jj.h�Д���H�0��BZR�QA��@qv�}g�K3B�,�v�)`]��������Y�yV�{�zOL� c��4����g�X��]��9!Q����- �+/�&q抠{���P��>��d ӓiD!��G9��sV�i�6 ��:��P�~	ż禄�k6�5⅛y_�?`�8�<ͪ6 (�i'��>V�j	�;�v��7a���j| QgGs"J�*l����τ�2�Bo�AJ�vI"�'�V��](+�4�(r�����lɑ?�����&�q�E�&O0�"��)9B~mq���d7L7� �c	-�wӐ�ׅ'k���zu=&TYR��f��i�!�� 7�P��׼�
cg����+@�Y���/cےi�!�B*�1~A��f䕾�?Px�9>#f�EY�����:עT0Z,�u��j�H���*�_t�<�����t0�ƛ����V}M���Fh��	Ï{u0�mkBr��⑰;M���=ւ���O�^�{�㻥�6��O�������W��3h��_��o�?i���@V2z����{��b~� ɽ��\aҔ�����>�qyd���O}u�C���n��y>�e�r����D-�u ��2V�55��~5U ���g]���<wnNu+N[���s�B$$kaq�5���4kCCQ�2} Y��9O3(�5���(v��r��|ƒ6ed�u[m�N���`x�dOs�t�O7h��O����FXG��%O3w�2�E���RV��	������yru�5J�-������>m�ĽQ&�1HtfOv:��$�fp�� ��SU�Kꀔ��g�_��팯_�_�3-��Ŵ�c�:
+�	ۺ��~�}�A���+�ц���S�}!j`�9ЉN�s4�7~�9�ƭ"���z �9}�[��i�{@R8H���iZt4u����r�|%��W�;7�}�5���S���k��E����Ǚ� ؗ������2� !����ަ@�mư�p����2	�%����V,��/�g���E@��K��ALi�
:%�`�P���M��O"�����D�ʮZ�B�W"mx\EH�H��2ʤ��ZS��G݉�?�� �j4���lv�ţwHg6��r��0՜41�F��i��m��̤[t� &��0��xêd���i_)��n�#�7<qe	�`QM��GIo���{).��D
��mø����m1�t��)�'p(�i_5~*��0�X�֮��P�y�z���+�?�X��4]K��i�\;�0k˃�MŒ\|b:�IZO� ��D��?�@ԡ�4��,بg�t�"P�ih�)�,��8Ic5e�zG�IO@�,�~�K��-a�8&n}��M���ůO�^������Z��7��b�e�Y&�����?���n����9��@@���\+)U�X���r/�M�Ř�>�Kg��oLoR{�0�v�|jս+�C��n�'t/wk{V�ܵ�ƎT,lﬖ�N�i��5�v���N��d�Jʤ�0�[~5��IU�b��IPr.� �ù �����WY��%�|�`7?�0E7w%I0��{�N�|�+zw�D��$��" ���x�ݸ� ڛ����X�T'ͻݣP�UOA[���W����ŀ"J������D=��V-�	�y"��+t�Pa�<r�"L�(��p���6��>��5Pzn]��W���Mg7XA�b�@44c�\K�G!Tp	�<�n{�Қ�w�3��XMfՏjΩ1&��JpO _E�>���d�z�K�[�6�$ɞ�ӄ�:|l
�3wۊOr c�ͮ.{ ��k�������VH�F?^�	�sa�F����,|�4Ѱ!�J%��G���[�~a��p
�V�?�"_ʴ�Z���4����{E��ϖX��n�&���*�[y����H�YUǌPX�`���n�����p ��xz��H��%XO��o[�����R`�[� I�Af|���H}�n4n�F�.�C�5�ٮ�jWE�}�8�.i��n|�,�O��OF]o��˙�$��|"�ӛz�?u��!��}"'4d�<�$ğٚ�d8�~�h�Z+�Ĥ̭������V@.��qE%T�ݡ�~js��f�J�e�dgl8�Н�^ �A���9���&'�gf|6��Dh���|A�j�mȩ@Whq�Q�bjI��t��<5���_�����g9Vl��V]�fyUg,xx_��	���w������d�Pb0�+M�Ǌ��>��.w]]̹��p!m��\���!$�v��Iѻ&�q;2[3�v��.���яrKE1/Y����,ַ�z��t5N1!G�u�`E�`��,�%��y��Ad�K�hn4]��XR�U�����1�/�oF���5��Ss���,�~y��oP͓�&�^�5��9Y�/����@�NN!i�o�=��S����!���i��b��kq|�7�����w��|Es�
�T���:&��f�Jڇ������?���9RhʾV2t\���*� v9eD��lԽә��Qn�2��+�ﵾ^@�_�(}���X�jɅ�`GO�ߠ#��'�>0:7��F�l�����Tb�<ۥm"�=1�UG������=֖0ъ��ٞ�OZ#K0A���˼-]�����_�N�r�ՠt-Uq��~^@�HK�2S�U#��[	��N���
�ݣ�az�t$�K���@��(.�B���F��{���/Iu�E}L}0킆o��È_Ln�LO�]�MM5#D��2��Ӑ����Q�n�x$�ע!�s��@7���w��92�d�JR/�w�|PS�|���~*��3Q!v����r:/FDEQ���w����A(�n`��a.��LX�H�>kF���8ѩ�u'��>X��aI}���T|m��n��h���p2����J# �(Cd�������y%�}Ę[��j��������\-좛B�K����r?%���&NO�)v���6�ˈH�z��ۉ��>���3�}��IGzP��[�C�O|��s�czæY�4γk��pzƒ-��	A�z�|�,ᇠn_<@�vP�Ȕ]��v(@.�������q�D`�w�	c�<=8۲��-N��%ߺM�I�k���:M��s�v���&��@M}���?jj�#<�R,���s����YF��T#�ê��!���VE��f��zb���N���n���lȭ���vj��Ch�.)4�Hǅ��͂����L��g{ڻD�b����_�7��.������!7l]�І�x�/��Ҡ�+G�}L^a^���2&���y�9@Bc���Ҁ���W�R�E��
��S��6K��DA�Z�^*�dj׾4�+G�)��ϑ`�,����&���l��h�RZ�����!��J��Ǥ�F��eӕ	dE�R�d���3�_�P����"�$����c��D�6�k`��{:2CQv�p^�S3��,���Y�Z�h��2˩K]�482�cX��N]�X��C�ήú��x�X�P6橾aa�	P��	*+�OFX�P��?[��F��Vr�&�
~��>J8��/�?d���1�[�_����?���@�ў�:ʯ}��<��O�����@��8�m���z?{�?X�na�Ɲ��1�N1I����,ep���e�0�="������.�`����4!s����j��@3�0�G	�����/�j�Q�Yady��Y�[���Xb h95�{^�lGىk �[�R�>j��[�7��F�8�ǭu�l
��3bz�'�����}w6��f�a���>逈�<���":�f>�3�R!�����t^�x���"���u��2��<������2MZ��?�Y�5<��Z�%�񶹚�ہ��3Q�}���tIR F�~�3��K�m�ʒ��n����r�DS5����K��7d�%^ck?�
XM� �<��Ԭ[�M�I�y��P�ۄ����7m�,�}"|Q��}]R
�&��\�iy��<A���4�kЮ ����4�Θ�����d%Lv�:F}lW(w�fa��	�a�<LD�*�?���v��2D�@�L���X��H�Xg�ߤ����Pw%�S�w�g��*H��^�@��㗡����m2G��{�d;w��[�Z�`~�I��Z��G6]��Ef��F��
�����X)7��ꍅ2|��r㸐>j�Ӌ�������TM~س) K�Zԯ�Pq���I��"7g���A�> 2�M�g��2ITŨ���L���WY�N
A�z�b�	Kc9�Ha�_3�&T��l��k�u�nV=1@��l�>3�:?�"�W�T�jǄ- /�	�<�������j�%~�����c�:1ٍ��	E��Æ�%��p�g�q��h!�4��P�KT&'�{C�.[ba^� ��I���c��8��<�5+�wv�g����W� x<ԏ�ΗO|�8�{3v�M�pExT��_�R0e��nrѲ�r����:��TL.������See3*���[��<k�<���(���֧�-~2�j,�'U�gr����X�+E������g=0��]c?,��]{�`gFp!Bw̦�Wu2��QW�����u��-�FqC��w�O���Q.��׀��6nY�+� �K�ۯ"VO�{��FrJ��ږ.��)��V���� _s��"���D6��2x��y4w.�~琰̱K����!oi��a-��G:ֆ^�X�P�;�4����q�3\�W�5�b�7�ͪ�.���pt�)^�J�!Y���uG�n�\?ˑ��5Tq���B�$�����`��=���"����U�8.��g�K(@�*Yh%u��u�34�֞n��kl������ee�(���-��d��x��v5��#Q;�����&��'d���H5���v����?��ablrS������_[�Y�<���RT��J��$����vF�i��akL��2��T��f�P�y+Mkdz1�X�s�D�e/��@u�E+��˝��h��l��H�w^��:>L붠bDf�qu�%e�<
�T���%����p�E囿�*�$��i�9���#'���aK�_����3�w�ֽQtZ.��#p���ҌS8s��M?>����J���Y���R���`��BM��B(=�*��4ģ\n�4 �X� �)�1c[gJ���-� �f�Z(�����	��	y:�Bdrr��Ҥ|���wL ���q���fSLv,]>��o�z�[oC+���ŕC@#�^�n��p�s�홪R��<j��!����j�0�����j���\XR�\v��Vd�~�>�0q9'���o�˴����O�V(r��,[k�iִ��.�T���xE[�ӸtR.��L�YĖ3����)^K���&g�n#V/=����3��q��vaD<�����r�b��c�z�k%w�g���G�َL���X̜y ����*??���? �.�y�$�C�d����ڽ	��,�7���j��5�3oWTQo�4Y�$�U��ACn��7#L�꽍��0=v2��ݹF�#�.�ͮ������\��b��`6�]����_�$�Ke�4�Z�ꖘ�rHn���2A�|�R_��5��Ι�9"�d<�X�����9�� 2`���B���_�
����ϑf
.���߿w_@�y�s_��T�Vxѫ�t���V��!Q��	N�x/W�$���7 �̡���E8�x��,�-����5-ꮹwK'{�4���%�:}$���-M�%\�w �(�x$dh9w*'Y7��r��_ԭ>�t�]E��u=�D#���T�˭",���c�,��iRV<a�O�i�؈�D����t����{� �\��P��_���n�����m9��	MCixR����	:��>���f�.K�v�A�y:���2�rć)ӅyɏQ>���0�b�=B���dԠS��̄� 4%�y+��y��L�{��1���B$��X]�0�bP�H]D��I�{�>���U��
������r";w��:0z7M�A `��oBf��
��3���v(V�2.�__9�ģ�\�a�p,Fe&��]��P�,v~�P=���9�c�I�)[w���k[)a�/V�g�G5�����:��e�͖��H�D>Oy��.��\S7��d��B��Y��i�s�@U���)��kLr�߇�˜Y��.�^���߀^�ea����n�VE������.��ԭ�xq+[��d�i7��u�qe�Y�s8�$��:�m�T ��F%y,+�k��
�~w�^q��3�e{6
WJ��%���R�I�Mg�:B;�Jés�V��LD���C$P�>�@N��L��Y�r��s�ݢ�p� ����tŮ1/u�ج"߉ߛ�߬��z%�|�h43��	�T[0y��r�=�D/2Ѩ�G�L���	ư������
�*��0�I��n�������>T��v�*Ӌ���mp���nwi�:���I�0�� DF4�Eȳ,2��ӄDjo)������8��L�-60/�J8m��w�z�m5 ��s�X��&�ylڞw̞�uey�
�F�H��[$�@=��!hT�v����g��o�B��p������P��xz/ru�a���F*�uo�*�:���b�g��p���^C�i��sx��Yg��Ҙ����ӳ�b�qI���5y�iF9�����ߊ���r*x�:�T�Gծ�l�t o�Mw��ܨ�j��7�s�G�IF.�����ʂA��4���|�-b����[ꃅ�-r]sf(�(Af~=�� j}�wNz� �VI][��E�I�'�(��|��z��2|�I�8 -I-���A�t�q@�h,�G�@�S�������(�?�cW��r��׮��a����{i��ӝ�8l�S) ��hdˊU���6���M�$��q�QS�w��LbD��q�.����G��C89�<����S�7�1Z;�?�wC׮�@��3�W@�m��ӈ-b�B�qBBG�l#H;JFe��eU�:�l�^�f�&��,]��t�W�����G�ك�7�8x���Б%rg.C׋�*����e��mP���*��.��hw��=@B�WM	7��%�m�l��Aҧ����0~�#�f�Z����;�}IGE�iS=@������
�����>{�Q0R���0z�;�b�E�R!�]E�7G�1y��$2�,T��D�$dP�)�-DE�rE�B&g�6P�����f��axPZ�&.m��=Z%��AO.�l�_���DMj�u�6���W-T�e��B��\��<�>x�&�.�ܜlIF@�&C�R�=�a�u�eejjzN���	����_����]��Ȩ6?�iB�)S2��+�����re�� �֣(�Ƕf�w"%��?wn��@�]�X?���{5}_���K�jB�'���;*��6��z��k'���7��+_c?�L�r4��"IHz6�X���H���@p#]�O<Cĩ�A��R�)�G?�1גbBÆHV++m��<H�	Lw�{�<�SQ��c�l�A���/�����Ǽ��rd��������o�ڈ��ݺ!o\�~g�\S?l�ؾU �]Li�z[��l�4����E��4,v������}��83>1��@J
�p�B�`���⥄���.h4~�e���/�5�� �}��]vv����9�`7���>8�tNҠb��9u�-�5��]�_;P-G�g�d�g�(��Uw����Q �I�^�xx8�Ar�<d�E�H��ױ|�D�T��Yjn7����}*E�G��0N-��ۯ� a_A��q�xuAP6�+���Q�%t]���,\������,�� #�|c���_�w�=H��[�7��;�����Yfk-z=��$<�s�'��KUF��e3�G��e�[I��5�WS��ʡ�����g8/�"����u��WQ��T��=�3l%J5�pԓ��=�,��Y��l��{i){�g���Cn@��;�Һ�<�Mɗ��k�{�Ր3pS.��T�ڻ<��g0�Hq���u��b6f�2i�R,��� �t=�.ڰ�����*aj
y�&z0~���U8�t�A�5q� ��/���(dݹ�z�@E �?���W����@���g��WFi.l�Q;H� ���o<Jϥ\�r�QkP꿻���hU��3�?K��)�8{lqx�%�n�z��^�i���C�9���?�
و�iC��S��5��p��Y��	��,(��s�:��qf+Ry���$�+s�o%U��ltH��� ��OG�)#���Ӿ7����^i-�Ɋo�a�\\��/YEy���PpA'�w���6��,b��8��!�M�˾�}����]<�
#!�D���Dz/��7ܜ;I�9Ho@���ƳL�>� kaV��1 ŀ�4�4���B��V��VA��>�)�������"����}�|�3p���s�A����H
�m�مu�㗁h�=�0�;PusH���aC����;5��z�g��U�'K��i/��-�a�*dY��I���f�Ѝ��'j��a@&:b�*8B2?z��9##�Q�D�V'w��zjy6��c�./�[Vꦆ��L*�z�I��GE�+�␍{�gY_��E4�E]CN�LlZ�iΉ]�84��{!�L�p��(����ԭ�H�(��՝@�d�q;����褞�"�HdQ$|�ڛN�'�����u�՗8#ԇ6ϲ1���-�AEuu��&��d��)UW�'S��a�Wȩ��ό�SN�ՈD��ͫ�z�a��=�{�7�>�B������}7�R�pcqg��?B�1vA�@6����-�p:�TCl;�u��t�(uﵕ2��	`nR[���/ǚ���֭���[h�mϣ�`���bz+���VĂ[�Մ��=�P�k�I�-׌� <9�������2�#c ����cҷ�?>�T�|��u�Q�ǋ��v{���-�xZ�����0 =��<�kV��DP����}+܆��+�)�D���@D�J�o�R�R`�{n\{r'��6�8��g8"�X�>�D�]Z����b�Lɲ�`ѹ _��o��P�a0�v�����q�Q��
�Il�u�aF��N�v���G��J��)U$�g��������J4Ҏa�DF���fe�)5���j:�99��Os�e3���ж�X�"��\�o���TU�\0����>��v��=�uC�q�q�M"A��1�i=�-0p�
Rfw|�Cd8Pz�	;��q�i7�s�9�KH~+�����Gw($��X/��
 ��sMa}Qfs���[flH����e���	-g�@��\`԰�!�$��0�jB�W�������U���u�{L�/e�tw����4c�j W���}���Pӈ�+�J��<l��������F^&3�0l5�� �U�BgjTLD�6;�Fu������%Ց�!_��Ǘ<��}֐żI��g��Aۮ]�P�D�_��y��$��Q���Ŏ�Z�w��{/gl�`k�('�:�rKJ�v�p�'B�}k�*+�J��B,k�i��,T�Q�S|��z�ʱ��	����q��{v��c��W�t�[��r�'�'�%�S�oj�O��w�6�?������z�v�򥈣��"�X�Ұ�nֻ��48�t,�L-��e-�2(Mt�,�G�l|r�sX5�˳/�v�,�'�ʬ]?�T:{�7���H�	L�=�X�j��!�S/����eD0�L�u���h���tݑ��T�~�����{#刜N�(�I�`�>Ϭs:Zc:���w�����+����d���7<���_t"�HE�P��O�]�X��3��B�祗�+�ә0Cm�䫴����]Ej<J��U"��n�_!a�\�Їv����>?ĺz|��J*���08ٵ>�A�YQ;J�Y��@��a:[�`�i�G�B���z�z�������!n$�j����:S�E \���f��z��S���9G�J`�1ق$V��a�/�_��"ħb��B%�����x2�vl!�Nl��C ���f����B�� '����)�����8�[FR��\:!�����D�C��_�j���!����p��h,�1
td��V!X.��p�m���|��h4r0w#s�N!��txi��G�?d-�����VN`>NJ�U]�1M�e�.'w��a	f{i�0��JK� i� K�ƪ�]]��f*M_@��47���7�	�*1�+1C�[)9�5e��@�)�(+ �.�3��!.��}�3�C��rW)"��x'.ֶ��!�|1�6D��f�pk��7�I�Jqe O��>,��²V��q;�9���|���Yh�hj�<ß�IX�q��ga:G�Y�fFo�J�!!hJ/X׬�@g�Q�^�KW	��U0v W���"�a�ҳ�I�>�x�����l-�C�u14�{an��\��B`�p�������Q<�Z�ɩ�629��Oݰ��4!�D|�rN$�/*������Hn
��f��7=��?��9�B":zj���	�N>U�oM+�]�)����C �]+F�p�u���wR̸�;�E�<�E?x[FE+��  <b4� �״O<�]�Z����~��.�f�^9uPL��W��u��G��̧W�};��$R*#���:�hLĞ��ﻞU1ӉX��;�.@/v����$_c%`[0��u6b{��$� �I,i���n6����P���%�������I/��v?K�@��X=�n�g`��ՃV-�+���˪����ʲWJV��C�:�a햡�E}����^�#X!�Y��k7uD�p���� K��چ�E�kI��vR"Y����R(O�c��:�U��_�&5��/zh��j|1'`���>�T,�G��1�׸����rxvY�;����L`�_0�V[ġ�:ܚZ�۔��X��M��� e���U�M��3~�F�m���(A�5�F. ��)�@]�#�%������Z����~�Q͕������I��E�h��Y�i�w99*��~w�а
�d.��l݋�x���hd[���"f�=�n��������qg�	��]���P(ذJ�7)^=p�f"봂^<:��P��&~��wp�,�8Hί��F
\P�5Z�]��Q6e4.�_FW�,�����n�Z�]3���6�c��4��[�k��N��i� ��"P���Q#k�l�o*x�����O/�V dܞ�LRʋ̕�|�'D�@ۥ�	7V���Fc>h��*ƀ�̔�$YpRp��p�u���Nz����Z�Z�l���{���4raXoa���`�O�~��o,����c�����	�ׁ�>j��7� '�T�$Ma���2.85r��u�=� :͠Ůg��M.
��Lf{G6�"� �0��r�&1 T�R�؇Q�Q�BB�C�|ٌI^g�V�ǁ��]���/b�Գv�m��}�t��r��`ٲ$������C�˫�س����gu�+a����-�R�\���D�tA3հxL�C=�z[��>�cҹh]q��݊���|�U���Jf'O�eUlI��&w�w�h�	��x���mC'}�<E�I���2����y`�؈x>��=�0������O�(���h�� 	S�EUX��+l�b�a�d���l(�.y���d��vy���+vB�-O�o
�X�� ��k��cB2���58)�q$!@�D�\�F`~&�$YT�p�^Xnt�'�_
�#��o�۪��$�{���8�NG8�\�?�����5��&N����0�9	��όٵ v�_�����ԌK�|�
��B{"J�Sw�vO̿ԉ��3���v�-�;���Bi~���*;4FM��%Q�<#���F�;:8�$�l�d�:�Mo"ibJ�O�H8�^0q�R1L��6;��mE�SxJ���[}zB���$6 }���k��"�0�zx��@��c��G�rAs��j�4I�rN\�T��������_bM͏��@Rv; �.�?���S�MtP�= I�ţ�K�C�(��?iyÍ)�z��A�$G�ǈ���������{�>r������Q�X۔�7�UlQC�`�ת�A��<$��88,������þU�������WæG8���x	j�Ұ׷M��"U�D�0��}�?���d0L�tξ����gww��1�(�e��a�~H�h�қ��]�H&��M҅�L��nm�^M�WnS��C7�'J�{ �Y'D�"P?+jxa4u�Vɫ��Ŕ[��Mfܻ�g Ms$�5Z��
lYu?�`Q`�Ѫ����:��ű�ۿ5F��Uxڣ���0���'��7�Zǥ;��+���|���{�ר/D�[�N,tr���-�����6��ozL�U8�[3��HJ�{���l# b	SCP��.�^���2����ˢ�ޝ�ȯ"-�5#�BF�eaN�����>,h���y��uVvrˢcԅ�@�QڮVlsh^�e��g\��[�1<쭚�B�%��cP><��ٴp��a�&�*J�R������4p�r���'���7��a�@�̊f�|�ا���Ϊ������<#`nK���
�
��M��SH�"8\|�I�[fha�i�P"ܰ�/���qh|�Ll��>�>�.��ږ<6��nMI�Ł	J�9�εM���D}��oONW���ቡ/]��i���u�Ĭ�m��C���5� h:$��+����1����_BO�EB��S׾�i�v(aU�5�R����~�/ˢC��Z���+k&{zt���F_��YxPy�7ѯ;# ��>%DΝ�k;�,
p&���q�9p��mħ�x�R&xY*.GJ�U�fF�~Y��찳\q���F-M{�r���D1����9�����ֶ�x�'i���]�roYn�(���+��$�M{��RA����>	h��W�9B��;��ī�����!��
��RY^'���^׈2DŒ]����� ���E ğ�S�}t���K�n�p�|��q�[��d�E�r]�R@�?�1�Em��+`fSJ�؊�tj�p7y�Ǝ�Հ;�E��A`*��t��ٮ��`�{��m��������Y���b+��h���a��m�.��}SQ!z�r}����d)�DA�
�I��O����ʉ�o�w�h M�BoY)G|�>����*�%���z\�?��k�	�?S� �m�u7���?�����]��*�E�"�\��3�J3��
�l=̼w�I5X'֙i7Q���˖��q ��x�BM'�NJ����͇a4��10���C�}��X}���rIK�>���tf�i���lu �:_ 'K�mhl*L�A��J}�͎X��}��w��f�#��q�M��YM�G�*"��w_������m炟 Ay?��F�#��VF�66�鎴QW�Գp��f` �ڹ�>;a}}f���̋����	y����szA�[�^yu=|y�b/孝�|��a��K[(�5���@i����X�d�:P�d���g��B�=�xfM�zxiO����]\R�8FC�+���m �.)4b�������`��/-�x�����f�Jڟd(G�;B0��ͦ#.5���V|qG>&xP�m�J��GXyF@! �۽|��j���!�Eő#T��<�z�s��g��C��`�w���꾎᭲*���ïd2�b�84E_��I����s��\�8�1$����1sv�h;��6d!Y��R��O�z.6$g�Q��	�rl�����u[	������q�$j��	�-o�ˈ��VJs��r�D	��FO��I��)�@�o��*+���j�t�͘�/�,d�o'$Zղ�wT#�&= �oq �۱��鉁<
CI�	(��b��%:/S�3r?9Qmw�hŝ�=�7Gs���B�_d+�( ֒n��gVS:LKp-�Sp��������Ա���z>��=AT�8�q���`7eKk����#ֲ-��ZB5��7��M���Wrd�雇l�G'����̔����Q$@
���Á��6$E�I"����w'xV�J�g,X%�)c�}�󞱩a 3��1�F�qE�Gط�O�#��V7]J�R
�$����H��o�ŧ��/H��8���q�%��^Mb�Ȕ(���ΐ�^�XUY�O���j�9.:�+���~�,͜�ؾ�c��C�F:"'����{����b`8�@�h��=���&�,'-�3�����yo��Q�j�o��Y�Y���濯�ݬ%G"N�bL{0j8�H�����Ze�}?V�%��||A����g�S���	J�z{��V��"��kv7T��acR�p-U��re������γ����l������u��;���VYC՛��ۊ���+���|��Q齯�(TiA��Q���Y+�
�Ey���&p�m��}�[��F̨>^'����r,�..*��^�����1��a��l����'���KRY�C{���,�}���n���N��?v��?�@���L+� u�dp��m��w�����45$��P��}� �������.`k��c��pHk>N�0IR7�U�rD9cW�/Ace�d��5���RGٓwWJ�gA�ڠJ	�:]r]�z'����*e��a���=��5�?>%jhz�Бћ�xk$�Q��G��7E(�۹�;՗�w%N��g��|��XD5�5\���Ȅ�U 4W��l�	&�>�'(����J��K'UGn����C��et����_�_���6�@a�9ÅRM�Ki ���$r-}���q)֩c�K����{�%A�l�9�+��.�)�|��.�1+�
#�>���0o�u�G^84��Rv����k,oUץT�\�`wEBn��E��k�̳��2M�asŹU7���6Ե9�!	��@�1�ε3ex|�LAB]��1X�c��eg�R ��Q�*w� �p���Ȭk��W��o>$/��`�Q4~1@�zdxў^Ƀ/�d���V$��-4үQ��ُ"H�{{{����l��,Q����`Q�ͦA,�#�i.�0���'�!��ȴ"-hO�,�z��+9�����3� u#�eJ�?='yD&2�7�w���q�"�@�
i� �yn�㺸���g=�s�cj�XZ��ȇ6�)�W�
��<�*<G� �)�h�$>���\��q����J=����]g�_�:���"��K����٤;9*�D.���x�!��swh��K�MRh; ]�}	%R�m�{�B!P�~&h�\�cm�oe2��ky�<ԗkx�k���\��������~�6� �.��0�7���.�����	ř�޼O�	�?Ż'LRw����B��Jp��/�D�o�
d��1��j?zRTFQo�B����RY=�#CC}{BB	� b�˵��'Q#�i��f���VI��q)@�}��`?�ɱ%������i�s�--���-m���6��^��N9�A+��~�n���Ƒ��}0�i3O^5A-���qD�K�����Y{�tg�}�ma����YJQ�A��)�f�N�����N'j��������Z�"�"��$'6�KFD�^���|�a�\s�F{�j�/�(�ԁ�1���r�@��+:\����@����D֦�����Oΐ�x�`�깈|��5m�';��@�F��P+J{�=���f��ˈ�mX���3s��}h�ڏ�:�N�'�2F�Y�!:�a�Z�Y��8&�����VP�kr�
�{_\�)��)�f�)�f6g&�}�=�§�B7ԗ\|�KA�q���;ײ%�M�=Ԙ����ܙ��ڲ1�f���p�D,l:~$�4�Q0�X	��q�4�gۄ�.�ɝ��F�o�Hޤ�Y"H���U����b�)�D5�ŏ$���~��,?v`H��g�E\~�1���M=�@��'ؒQ}�,�*f��DT�T��Q�m���N0lY�V)B{�$X������(/�s������Xvk�����0�(��e%(��Y'�ؓ�= ��A�3r���q_/s�`��N{��1���٥��Q��|;��A�]3{�`M�n)�w��U�s�Z�O5�|�W�k�6��0�f�:��JC�k��@������!N�^��E� ��x��9id��)�j�b?$�D�md�1�q���%���w��TK!i��~�Yz�aDҬ�π��M�aċȰR']k$�@��T暬�jsgb�V�<1�d[ϹYL/�Y�[�Im����{�8F7�y��9`�bo�����qXK����d�ZlC��Q��m	�sS��o��`��܅���:��D��カ6(!�����ˎF�aQ�s_��P�e���ƪ��=5�8�8�v�c����X���yw汌o-�G��U���~ޖXQWn����v��mT��B����c�N�������K�/�y���]�r�n�=�R{��Y@��Fۥ�S����e�]X`#~)��]�?��m��]��C��V��O}�	�"���,�zQxPfW!����O:�>f��e.7���WC�ݔ���Qz"�4�:��u��wl�R��ojF[��S���,��N�k��E���h_Ƅ ;S��uY�|Y�to�@Dl���P���b�퉤i>3���+�}eԔ�e0���'5�Y�����st��mfh�w�{�)3K�Z�1>��y"���I�:0�����EK�Z����Y:�sީe�B��G�y���6'�Ӎ��ˇ>�Z�8B�7�d���F[�c�c����a7��}Cܹ�)([[��X�����Ig��w���2�Ў�����,�V���+��y���Zc����J3һ�3B�t�bo����	| sK�b)��(�ZH�����6A���f�#��-�z�eɯ�ɺAJڰ��	l޺��1FY�X,�З�GX �xN�g���KL+��]�����8�NH��.�SP�X�w��6���[�!��f�{ ��M���R�Z�!�����O�N6��v��z�N�t�ږ�?��,���K��=ʣ+1d�7�6!��3�� ףf^\�����G%��
8���ڱX\�!1�\,t���Jϝ$�YA6%g9��RF�4�Tw�u�����c�x�8Ө��;�R�}��۽7C+t��x*�&G�_�w��h�F�t�!��?�8�s��!M�Y��苮;3`'+P�;I�i�n�Q��$�٩�b���Q��.�+S�%��Ǜ����h2�~Ɯq()�$%��J��C!����h;r��$�<�
[�B> �K[���S9���Q��vO���K�����J�/�PhX��6��`�pD9��sk����\,���p��,UP� �:^*�T1I��6����&�-H~>��4Ԕ����@��}��ڈ�Q.��'�M�=���e�"��/_�ew ^TE.�4�«�.0C���B�K}6[�F[m��(�C=t�b���]i�.� �r&(>?v�CK-�k�2ߩ�g�?����?����j��6:�=^�W�Sݪ�p��&~�FL�{�QBv2%m������*�O����g���o�q��E����5N�jl��RO���>>1�Y-��/[���ł�v/�/�	>R�b(�jQ����4��h��i4�-����lub��I��?���s"+���?���4A�0�������A��5>^.�S���W�燏�p�&TC��.��6!������IZw,�,�V	����:�KLF>�M�Y�#��9�~ބy��ZF����|�9�d��zDc�4��$Of�m��I"��A��h��O���T^��舘RrH�(�z�,�|��R������
��S7.�i"�k�m�z4�k��s��X���p<.U�,�Ñ�T�R2L��یr?��ޔ�N&�*_ZDx���}��P��k�yH@V^ݞ�E2F�Ni���~��cI~��X�!?b䯜{[nr����Rֱ�{�y���u��@;_��E Fm/O6�T��}��d@�_�!A�F����d�W�1$��}~��<j���E��=C�d�1�"���2�
tk�\DB�Z�G
0\�	5 <��#@�B�NR�7��p��I����{���屑��CD�4/�+/� ��7�Y�
�d�';1�j��Ml7��b{��momn4�}���?S�ݑ�i7~��8cb=�MM��sF�v�"O����ƀOo��H�R	��~��4�S+M	Vc#�!��zG�1A@߳��Xx,7=�qЇ���@��W�֙wp�9l�7�T	"��RL����57�B9T\"�����b�aH_����!5�YZ��=;T����>���? ���~����E�gJ�AIN���	�B�D�l�)�wVʣ(��#�͍s5�27J���+�XW�ۗ�	����(�� �:"���9��+o���p��
vo���������/�I4��QM=�� X~Ҙ�؁c�7ի�7��8�E�d���h�i�hS���W�%���ObړI>bv�w��N����~Q���&Kf �"'�S<D���}�ε`�(��R74���E]y� &W��>P�`�W��#$} @7&�H�:Zݦ�m4�g��3��%F1 �CVAQ�q(�T�{ͻW,4�1.�6T$H�Y��5"�[pYʉ�)n����4@�T�8���<�qQ���$<~��^x�'ꌰ*o���p���QN�dB����˦��^0ai,��z;���5��{6�����q��{��3���m�/����"tP�Ăm��߰=*�`�Ԉv�klb����r�;J� ���G]ȷ^[S������W`��]����O�{�"C�({��>���F�¢R��R��ɯ]۵
#�k`t9��K\u$(���+���b��ou������D�QT0~�����pq����5&KM�WyxQ����9���Ԏ#�Pv>���Ib~�'�i.��Dr������($[yR��/Y�@�wEL��EL��M�QUs���@�-)��h�%��cN�+����Akt�W5�q��'�P
3J�,�tt4�����1���� �������ݪ/�裂���������6޳cu068�Ej_^Ҡ�{X-&�;�=�	/H�匿�Sm�>p1Von&��!�:ۀ�iS%�f�� �~RNM:�?�X�{� �Q�����B?��=�=A��Dk�; ��JƑI����?��6�I�n�:�~�_$١���qT�q1P�B�����1C�	��ӫt����U
&�(sPUH_�|��'V��t	�%�@y��<�zIN-�c�*|���K��M>�^hX���|�i��E��<6r����#�UC1�� �,y 02r2BN!Z�M���sD���IW��
� UP�'�wԈ+��D���.$��,w#NI��D}{!�W�bh���l`�/!wN���������\P�W�T�@1n\��{T��n�`�ˏ���N>��p�V/fC蝝<�t��i
���l��e���[҇�i1|��c^�Tf���M���C�,k�к�ju�fc�J��:�^ڝ�
si��L+���7'���ʅ6��w�T*���aH4�93Yi��-�X�%�7iy�H����_�ч?��I&ME? �v��g��F�9,�l���(r���1�">�Ҳ���R�.�T�*&��bs-��kfIfH���w����p 3���m��ig��E�!9��8x��<��������9�y�D�w�O	2�`�����Qm�F�5��w���Ҥ��N�c��?"�f�p��S���n)�W�S3U������ ��WA��׿��j�!�Y ��9#�i.�jlLssb	K���c�����
B40��@q��F�DJ�D'X��`�\阆��.~Bj)�M�E���>S����6�3���j���b�cO!���{�mrx���ɵ�[U�Ur��\���}�-�J�j{C~��q>����J�>���w/U�m���I�j|��lH�5_z��� �'Q���AMٮj{���D�|��I�=Sw�W��?��}L�����vP�Y�>*P�rQ�z�N gI6_is�JK�T�5V�qC��I��f��lϻۂ$�2�go�j��U����G��N����Э1_%Բ��$;6����B�I~���}a��`:~�����Y4�<��=�㑳��V(-0Z`F"#��L�XL�m�}�v���i�9K���f��`��{����r�$Y9yy�EG�W�� �ǖ2��Z����WSv>���;�Z�G����(1��5�2W���})�&����fJ��՘y�4j*) h�D��n�ˑ�$_�^�1��v��,����)��b�JZ��Q��$F���,.��5�2n�G��agH�Tj�<����09�A�1�[a8�S��ڶa��:ϐY��z'�ݩ�|x�GT�w8x�����W{MKl_���d���k-?�D�oM��,@>��L�9�[[e�
R�p}����W���K���WJU����s�z�9�X"i������1-��*��k7זN)��a*��@k��lPM ���X}�g���X*v����y+�P��F�̡�|�Rs��h2~�1��g�kl�[Y��j�D��<~p���5�1w��a�J#�0�4�h�E�z$�?؋Wc!���W�QɌ�(�f��m�԰�?��_��=�� wѿ����*���	���@!�jr��+=f.M�h����ŅƠt�;�y�����֗�d7�ǖ�aüX���K�T��;���֎!x\|�i�F� {1'����q5�3	R�H�Mn�>J��7�˜+M��P�b�4��^vF$%5�9!�Y�K��~����"3~���A{�g�s��J�賶�M;���Z��I`���*�VKF�- �ڃ�]e�_��u�ǭ5�L,xŚ�>� :}����l��m�]Ž��~ ���Z�����[P�`,3��U2@nZWI84�?cL��E�Q`@�Q@ �np3���4��FbC�Ef��;B[c�!�un���j�}�*WP�ɰ�V�N��I�������6�$��U��f�.�u�&p��>�`��B�������C�6`T�ԏb�$ƞ0���� tf�������Twq�ʷ�|�m�V��ӯ�C� �C���>4�IO	���e�iU:[�mo�������:/$~�r�	��#�
�5�8k��Lʙ�:���n|\
�;S)�5�7y�]	}k$ct"i\QĢ������C���4Zz��G�,����GU+��Z�J2yL���2B��ze`v3L(�KS��J<V=�D�(����u2���j�Ȧ�����s!d��ÃQ�f=���"K�k%]���Kw�bl$I�E.5�p��v�t���6�;"�c#�\��$����F�F1�X�4��0�rx��+�J2�c����5֕0?��'��ZY���ז��*�1��	ջ���C��m�	�O�,��ڔ�n��m7b����X�x�Ƿ��ԹE���z"���Mk���}�?�DOnn�; ��"&�[�d=�ߙS�����e���$���q�8<=�(=��s\ƕ�N��M�(^������y���.}:�n�z��5�2���c�I�j.�eM��Fg��A��Xr��:2 �khB�c�_Q*Ts4�I[G%�SG�p����i-�!t�����nT�VeX�~��#v� ��W˄�Z$����s떣 ?i )���,)��jq��� �E�-d���Kp���K��0��a<B��^�M�ڍ���$l"y���3�:ygVPE%e%2���ːYJ�7�R�zKkWYM|?�yl����G�Oy����\��Hy�j9��Z���4<�60�)�Sc������?���0z����y,�O%�_	H�OT��i:����ã� ���y�C4�~Z� t`��luOM��j�u��f�^�)}��  ��߀�����f���x��!;4��R ����`�;�j8�&:"���P�#���.U�K�uvmJ �V$����e��kdD��a���AJ�y �aa05���'<s{av���N�Й��6��ѰȵS���)�X�=���L x���$r�,?����o�n=��2�Ե�����0^��Ls�B�)�$4�L����������W7�j�/�sFi)��f���R���8��}>��BU�=����M������5����/�̍\l�&���֔����1VkL��
t�I�u1h�Kj@2" Qb���\���,��vC��tغ(O�YC�,�9��a�R����*B	�m�ɁtD�Md[݁�B)
-�5�J$�8@�b�Ҩ���Ò��k�!'ݡ�-�\��2� A-�Y�e� �tD�|�S���n�*��D�K�fTA,�8)�g-���|%<�M=�/pc�5�w�$�wD�yMP
�����DU��`)\��01a����%�C���1@��|a�5��|��稀<���
�[4�
���&�����;0���dR�K��JG>����b� =Q��{uh�lQ��d���A�ީ{�*�߫9��rX� 25'U���g��r�N
�˯Q[�HQ��wEh��=�۬�V;�y����#|��Թ0�V�>n3�ky�h"�D}t���7��V��w��Y�~H�Y��Λߤ!���"%����O_xn wp�}聶��Y���!{�S��pՖ�*�h�aЇo
S�C�O>�v��F�P���l{A���X�~U�}�Txa��6���p�==WGq�$�QW��7s��M���1�Ss���<�4O'�,�ER�A`�̶�e��z�5�3���ڷ��-q���#��ы��}s��
����>�3�T�4�`ŹuL>�">J�����ϩ91�88��9���#Հ����7mP����G���g�f���yJ�63���,4>�^�K����4]�n]�m��·r#QF��V#�(o5�a֨Z[�(O�,-�E�w���g4����/���Wd�v6$�O��	#U����D��暮��5��O����]���7�� �?�!�K��	��cLߑ�B����!�3�7.u2����4��Ǎ���oA�Z,���%�A�+��>����D����\[<rs&�<k��+V��Gi�Sk[�n���=&�]�&��6���v Sģ�ә��I/���w����߂��=�K����"ws(Df��[��F_��0_t����t0I�\��M�B�:)Ւ��>��	T ����Խ)����u�y��y-�����6��<��!|�V�B��ݬO��e"B+#a�b C%+Ɽ�,#�>� %�H2��!ޮ�4�Q�,��3�6|�'�	U�́&z������4ӟe'F�ZG����_����Dx.��b��9M �|˝�U�׀���廠��hZ�w$��HD� ���y�9TcF�&�� ��1"Ǖ?2�{��ȣ��h�V��WJ��庄K�
3;v���[�3���}/�;x�O`�q)��ԅ�4{�j�B���x����Яt9��q^u'+�h���!HI3�G��1��6�+{�C;��u�jM x�R����ȸ��L1}�^��"�<$NgO7�L2�1i�*-�T��������i\O�Ӎ����6����l�F��x>) "��f6Q����y�e���#�!���ujw�e�������@�-������ԡ����#�x%ԏ[���SBO�dz��P\5�.��aS#e�p
f�����,d�c�ms� Y���:*4�Y��o�t�V�2�cj�
F�γJ٥�K0��&+PS�P|���u�Q!"��9��
��#��1����:��� �Z� �5�(���5���]W#��4C�:gv�x�W�6)P�ڠ��]�c�9-���+���dAZ��ɩH����^� �˩�٢͊�'�O��$d=:=�Q�����H2�;���p�\��]� R� �د:��t�ϧ%�h]sD*��(��E�3;K�0 �(�R����3�7�2��y�(ƊKq�:�jU��8�-������R�'��T���
�;��ӛ+����#�#J�==*;.�6��۝#�W^�8�`0Β�J�j>�E�Mn��o�l}q�	�18ۏ���QA�Ѓs���$�l�.6/�`�$�T��Hby�8��"�K8G�dD�bg��3��#�w���Up�����8[��T�M�����)EL��p�
��
����G.��Y
��������Gr��)|1�S��#�*���(����0���Jz�~��h��v��q䉪���n�{8��1�<�1���R�l�B���dD}7������a�\���G(�y`ɽ��~�g�~���&)9ܼ�����I\iY�E B�)�c�0s����x~P�K(S���9�t�]6�B��n�;q�	�C�}'��+2�����gH�	k�7��K�4��Ӑԅ��G�+��
|÷�n�`�یg���-��.����c��uD�Uo�Y�4�KG�jfp�{�"r��0"_zL������>�x�2�OK��P��κ�S/��i!��A{9.�YU��Y�	�!�}RJ���7}�m��E�����%4���Sq/%������{O��2nHj�յ�
pԸ�٘ތ/�x��H�'6�w�z�8��2�S־��?��d��g�\���|�D�^�P$[��?6d�))h���;�_�#5Ū���K��ۘI�mdA-T�����3��@gi�q�J�u��	��Y�3̯Hv�iQ	6:�	pú��YB��{�Ά���1|ĬK��*�_�j��H��U�;8Zu~-������^ Q��������Kh�'j�|х&A!�8B��N=��*��O�h�pİ���;S�9����\FnJ�Saw��I'�M�R�d���2/���_:��E&�f����{xh�YW�״ѣ
�ތ��i~�.Mq��q�g@���n�v�����9dtW{�`Z3Xg�����M!��T�F���ܤ���@��L��9A��g�:�󧞙}��Pi�EobFBc�s`s��tp�8_�[�[w]	<Y������:��3�	���A��ۚcn������nZ��7飮��y�d�J 1���� ��c�b��w��NFs'J�ʳ�_*��Z�eKN�v��¯��ަB��H��va;�����ϧ�{{��%�A��p��n_(v�ƶ�6_r�NJǋ�A��W\��^q��qU(>��&!��5��A>އ���!���l�K�b���+A?=��6A2�iG۠���C4}�4K6NG�u,�z��G��t趯ş���m�u'��N?n#�����*Y����퇊ppU j��:�'r|����u��z0G֝�s�=��%O���]L�ޘ`#�6�"�?��	�F7��F_	�Hu�K�t���G� ���D�u�NL����CU��q��Ф��5)�Г�M��Z����e�P]��A��i���>y^e�EO��GYpD��m��9���2ׂ����z'�D��C��$�X�D�W�6�)�7t��l"��̅7���xqbT������~�8�)Ff�v�s��͗�����d*�b�Z;�آ�6U*ž(?&I�zp!�`A~*��JȘ�1�HX$y���ʺn[�^�m�l��^"���b�TE-k��Y�<�7�w37�<��V|���or�b�\��"o�zt���RA^����z+�m�B��#t3��M+�%:Ar�,t\2�������d��ӆ-�T%Hz�W����C�+�|d�/�߄;��2��QI����ч�f`��NT�с��#"V������:��^��=��Q�3RO81�j�;B�F�50\-��u�at4�w�u����ո���Z�2ON,UY(�(�_���L�̔�q!����1$���@�_-��Qv3?��KV%�21�̞��zH</��wvi�"�ƿ��e��\�pC9�w�O(�h���hXy�U��|�.�!EQ(င�Gϡ����Q`�!����(�v(
 ��D��"s��^���>���W�hmi&�C�����E�|k6��GK��{E9�����!����0C�3N�0
O0����%K����*R^�7�� ��������:î4���\���
v��
�R�Q����ʒ��}� K��<C�Y����[����F�Q��^	7B��3y�&��|Z�X
����H�
��D�I';��yM����L�/)CTy	Vt��R��H�����F?u<���G�p� A'l�䉏6N�vh����B�[�G�ж3���6���^Y+�Pa�Z?�A`�"'��yӌ��'��3o`�+��Bg���%c�ՂpM�7� �?6�B�s�����*Ջ�zZ͒O5�n�+�nY<�81-lU��z*��̈��t���(E�'������ ����煽�w��e4�i��ә��h�
��M=Mj��z��߳�M'Q�Q�8�!� ���R����C
,��]���׵*+�����v�#��o�98�l�t��k��f��`%�x%�s���H���/�|[V�孠�gA�z
�\��XO�����P|����0��&6y��}��ZR��Gж��b�C���<��5^~
z��`��*���i3�["���)C��u�"���tq�[k�a*mlZ�Q��	�LH����_Q�4Q�8���r�Ͱ�f:�♕�%�(,I⚍È�ɉ����Y]	�j�_(�
����az���+~���p���dT��S�NS*���vcᢖ��%F�ifT�J7��UD_��"�TNA�����K(��uo�y�����؋p���g3wl D��{xC=�߅�L�k��eU@F��).�DK�t��q�Ԕ��h[�8sk�/���(̓(af9�ʉ�Ae|�l��5T�~�Q����)l�e�֊�uz�҆p`�"Y��;��3ʥ��Q���'o�z���Iv ���1ԗBO�^����uX"3�˛փeB��E/\f&E�F��Bۨ8k��B�B�g$���ch�I����:��Z��9��Y��iRr�����c��ˍ3HqP�g+(��`i���vu������+��H g�Kg4ka�Ȏ]�t��.����ߌbi�r���л����c�����mi����1`�ys\,�yxl��:�k�
r��l�4��E_	׶dJ[cdݭI�/�'�d**}`RzJ��9EN�CQ{����9�g5�y�� [�GHF�Get�x�ɞ+:�s���*��������n�d�Áf�`������9��'ܓ��v����[��.d\� �w��fi-�)�˙��Q�]��@�h���� ��V�a�,q�
�JԷjb跧tNQ����ܤ�i)�f��1�}~۪d�o�̺��d�.i���\4G�a�!�%l.zـ(L����Ω&���ڹv�%�y�_�W�k�����1F�����ъ���ͼ.�
;�4��#��6�/��!Ǐ��E�T�6���4J(\~h��]
C&�1gY��!x�$�Ji�9/gH��vж����!3�%f ˴��T�"7Z��L�����T�Y;�K�T�X���~,��ylw���ݵ$:_K�����|�ҫ��y�I�qȆ�-Š-i��?1���Y�M����F:&�5�ҽ�c:�����x�r]\�ՋM`��0��/v�V67�dͳ~�kr#w�׳H�.�o�.R�L���jׇ�D8����B��N��!����)�-�V��0Ѵ�*K�{Ұ��F�=4���ǵ�T�A:�����J|:	�+�-���ur�g�����Jc�3�U��OW��v����n���
�f����>F�/%!y�z��|�ﻌ�yg���*4ڒ[t Dw�猂�,�<�CK�&|�_��V��9��yX�J'<�䄒�Z��1��@_k�M�����hlq�nʤ� ���w�L�x7��ϓ\I��滢h��8A3 ����(tK�Fp�yL��Ҷ&�/�m��T�I��>��&���<��8�-C�8SB��F"��=I���5�YE��[���s�Y�g��y�}��ҏtG����x�{��WުSM�����N�&*5B�g�Q���Whd�����v
����R��A��� ��2�}�K��1
ڐ�g�V[˪�C&s 8�h����j�M�c��҃ =$�]H�6�3`��)5=椸"���N��5�K(�������m��j�Y	�2�d$]����@+1;�����+;0�����1e�>+8 A�ECbs�V��U�2g45N�ÜF�����_�s��w�f��i�qg҆�Ἅ�D�l��خ��Ѽ���������i!kV�l�e߸+S�3�dr�¶H?�=�R�A�!d���T���Bck���`�ை��o�BoUu]�b���.Q`��s���SF0o
�d�Ç��.-�#���[S|v���*8$���u�_�Kg&�əF��\��q�G8�m^0����	,� O�.͐�>��+c+|��h.<�m�`�l4���ʐh��َ���'CM	y��&o�Ŭ���+g/��G���{�h��%jd��!iA�`�Y�-�?|���1Kx�/g\�]ң�X�Zҁv�(xCu��@MD\�/V=����KTu�\�-� >��$d/��nߚb�Z��Nzb�e����J�9V28�w\��A���[t��R�2G����׮s"״mZ_-��'����
 ���J}I��ڽ�&ʢ�Q��@��Z.�� kF�-r�w�r�/�ݑHP��PD�Hѵj���;�Ұ������9�7�)���-&A�D$�^�E6�$e�U0K�i�����!"���Ľy�)@�vf�n�"Gԟп���Ëq�W% BW�qQ�_��r�)��jv�ɜj��0�:�	6�*���m�/ⲇ���Dy���P��6ن��4��7�̑0a�@:ʶg5�b+2�+��k�s��:h������Y��/�����JXZN�]s���tH�r(���j3:�X��s]�l/�Ȁ��[��^G���D�݇Q���9�Y� �*=�B~:�/�֡������Ad ������itv��(�3`�D��ۺ���UqR�HM��8=�HI��_!����7�~)?�Y@��6u�!���1L��i�}�홍>�����D��Y=��L`K�i�YaR_QP��Ez��Р�{�@��4�
��6����j��T�*�?薱6V9��Bfe��~�z�0W�h���%G%�,۬M�*`a.�ۃ�؜<ɖ���YF�E�f��޼f!���a�И�R�#�H	�S"�w�c���`>2��<����n~0���f3#F��	*�P2�'+B�սx&��A�
7<�[�kq�ű�|dD #�$x�4�`��Y�[<��;��j#U�C�����;�4;�_����P�[��Lf�}�/��[�%���aV����Li.7��>+����j��W�ʽeW��H������f���XA̺R�4�(����k-����Og��Qф �OԠ����K���hK	Чv[b�ЏcuY�� �L<�i�V��L�Ԗ(���ԏ<K����`b1�4F���q`�z{�!��T�Z�B�Ң̹��{|�a���p:v�c�W��ɖÎ�t;*-���Q��^�tbw����r�����~ ��f�z�f�H��ai����a�,e
�����c�dz��n��]q�{��9|E"ǩ�����a�@w��(^�d�����q��U%�O���dt���$����cJ�_�)��n��x;a��8�ܨ*tф>��m0!�9h��m�D�����h�e�0�h_+c�C��X
�($_���ϲ��|�c���m�=����9��֜?Z�t�,7?��U�5���#uեac�FPn��]kr%����`K��.R��6t=?��-ڛ�u�0�͚@�wO"��oJ��>����,�,��8r�O��ƃp����5����;�0��	���֍-�uv38F��%�V'ո��r�5b>&_�j�e�� xg�U�up<�{�#�{���D����$���av�FON,���4��~:�>S�kE��e��v�X��p��	K�a!\�hq����dd:��1s ?����!��$垏�l*%^*�ZVk74�CZwyY�D�: �8:��Fy�����)%���}�Z���w�OB�a����f��z�:+�tC�aނh&���n��	�� )O�F��%Gk)�^��v9YIq�wW��ò��Ũ^<i)�%�d��=؞
cQ9�j,{C�G�8�������J��>�ի������@�Z�`��ii�xk���+;7g�@GGi�O)F��h�
`������B�F�Pz��gBg�WzVPa3[c�V�l m����պ�Zu&���M?���C�/,�q�92�%iH(r�tzO(��o@�q_�-�)�p^NS���:��Ҳ< i���G�W��}�Baa�/R�Z1�П��ݔ�YĄ�mp���Q%α�/)���h�5�n:���f���E�;�st2"�����A涳�t-�A�y����@�߻��U��	[�L�qUɝgG�	?53 ׿U�JW���S�ɛQC�S���=���%��T�2��S��Z�KJ9k��*����zw�@��F�"�<ƶ��n��m��	[iǺ(�݆j����� f�m(M8BS*�Ŏz�Ҍ%��ƕ�4E�]���jAk*��T��I�I�*RJyb,��6O��k)4�<(��}ָ���?l,(HYa6+r�F%]=(�S�dꌈۋ]ll�{��Q<+Z�<��8Y�b�$�B`��9Sh2��dn�;���m����N�1�Jk9��0̶3� ��weU����[H}>���]<�V��O����M����Ź%a��}���]��$l�r�s!uj�Y툍��1�C�]��*�܂�|sɅO��ܱ{ *��N��)�fh�.X����r����f7�Y�n�]x=Þ�_�|w�_����k@c7ǽUO���%���A���ӄ���)Ű:�Ra��J=;��jG�dڙǗeb��Jp�ٻ���O�}���h��=�b�����[7���)ق`�L�ɛ �
�5��؅��Dĭ�r,������w`���P����;63�p@�Sژ�L�v�ѲB+��[����n�K?�u�{�-��)b-V#C{A���G��>8�7�ZF�h��E��~Ѣ��KE���~/�a��j�s��Me݊�8c�CdD����ӯ����>��m����5$��
)qvgL/�;���Ǵ�K�#)]7v�BĂ��X�C��-c(��叇�����L�ה�&F��U�(����՛#~��Q:���z���Aa�k�d����Uu4~�5�����To����朸Ju�3[%�$��?r�_X������-���Y�T6�K[�����C�<P�"�)GJ���x��t�����9t$�y����b�h�N�&�UN������ˋ=ꑸ�J;r�[�9�*s���~�V����BS:�i���G�x�a���/a�
�~��!kN��}�Giw��- �� i[�Z�L}J �~����D�/�.T��wO���\��x��a,�J.��m���W�c��8-m�r��~&��ĉ��	�~ncc�ݺ_=X֯l��@��/�;Y���U�*���q	r��_����ɋHp���ZU2�=���n���\La�N�I�`4%(rz?���¶���=��Ap�{ڱ����'4f/ÄQú�&y�]����]eu��ՔPz� �&Ҵ��i�Db����S�CB9;?`�-,�%H\�B��$�J��[&�v�[k��5�H�'㤮ɻ,�c2b�u�B�&�HH/�CSV[�=
��J�70�Ȓi��k�j���j�Р�%ʌ1�s�$\`�{���a�E�X6�F-R:�����	o6�l��J�������S}���I��GlU��	?�ʄS4���
��Պ�6,�:��:���'�A�����4��zj��(�e_�Ĩy�J�񄚗�!/�$%��h�B�G��J����E�a��t�=��,k�O7CL�|�j����U���]�-��LdS��_<�#;BC�
1k{"h��)FI��<ѱ�<�Ǎ���֖ ��&� ��ꩇ�����g6� �:޺�/s3���>S<�f���|��֚���!l�����;_�]~�	��Ò�H��a~�6��pW���w���ė��<����� �"\��]�%���|PŲE��5�?�J��b���wYh�3�H�o>}F��Q	��}��>�S�۬2�-��"�r��8fTǹp���.�M��-�m�d��(�(3�1*w�^��RX���-�XnO�:P�:�i ��z���k���c��+�&��!yXؗ�`�1I�
F��p�����t��0LtN���ө#)e	k�#���L'�K�x�V�9�'��_!Bz_Ac>��>�8<�o���5���MQ��=�\��fݸN"Bc�1�Ӊ;IZ2�N�8�tc']��ECJTqԴ3�/1�Z�I�@�O��$�p������^��f�*�V�x�Q�m��Gh�'�K��>�	���%E��랖��U�u��%��|ʡ�{�^FS=�:o�7Lv�3����FJ��h�������
T�22� q@Ӥ�]Q-O�S=0<����*X�K�m��JZ��ο��\�'Jr����O���(��6�W�2
%��8
��6��BӬuQ�uR��Y�j-���3�� l��O=m�&��2����cn�J� 3
�i�`��*���H�RS$��{5��y���L�.��.מ��EI�M�o����2�̯渭�]B�1�����`d��Q����$�vHC�(\0��!<�f{yE.��;�=�c`��eJP"�m6���K
�5e�;!#�?Is@��ڶw,�?��K��$��,��Tz�ŁzX�s}��/��ww<"W��o�u���������z�b b�L�ٸPk���M�]�͵ڶ^�r���&	Gz&�ŭnO��T(?]���O,��Ol���%�u{��sn+�~�{�w�7 ����Fd�ohS�CE��y�q�zsW'>���$t���!�ߓ���)\4u��1���e$�:�z�g؈&���$��~�<�!��v|�OJp�*Z[��>�*��ޤmJ��Z�ɛv���\�6����葕�38A��Ĥx@��sgt�lᘆ�	����Q2��Pֳ��W�!�s���HRMs�_#���sӫ�����G֭_�<vE�;��l���ٌ�l�}�ѫ"�(*W%t�-E�P�C��e�m��r���}q�Pm���PP�#�Y4ݮC�:�I��C��t�B�C�f�ʫ�J��3����Z�������� z����1qK0��u����ɘjէk����G7ڙD�P��'Z�c�>�?X)��*0ŵ�+5J����˺�}��ۑ��K��3���@�ۦ����LԄ;_�<%��(�z�X�Q�[��8cg��~y9Qn^$T\ύT��%
)�Ү�A� !��
���#}�x�صW�� ��r��%[��H����Mﭢ+͆�'�%<z?4J�&�:�fK<����S	ؖ �Y�o0�������M��a#L+_ySx���๪����>�ߚ�Q�]7˼K#06OP*���܋ ҍb 4�F�Z 0 '�;�F
�L����'F�;�l�?h�Ȓ�NGwF�X;2��$Ƃc�h|���𛪚�-��|�Vj"�H}��YeI�\��_� �E�P���÷A	$'>B���5s��Dh������5﯂}"|=�[k$��EX��Ϥ���\ђţ3�o�F����gWbxf���N�-~�h�;�7y宸47�S}B�C����Y,}�x[
�]�,�h
k��$�6?�~��V���Ւ���n�� �ry�l�$��bd�thՏ
)r���=�^!��#[Ua� =��AeO�f�'����oK�6�l+�J LJFe�H
q�֛���C�X��'<�Q�p]�^�|��<e�S.����fd�]k!&�
�I����b�wüvoԡK��d�_&
��R�������ЪD%_���#C$�=ٙ/w_�_"�6�����*�lJ��E/`�s�h�Y���J��v+n$i�ﯱ︇�h�N��L�ކ��2¨ȅ�p�1�RE���u�(&k�niLc�X$������Uw\4�U� XT$p�:WQ��F}a:�[<+����8!��s��P{� O\�d$�G}G!�{V(�N�7Dµ0�S��CX���b��M�h�ܓ�RR�~5ÜK���{ 01K�gTU(��I��C��3\v�%u��
��!C�`7(�9M��_�0u��Z�=�(S�U��o1����X2V�h����'�8��q�UD����w�!��/S���+�eA�[x֪?D�뵞v_�k�c��G�rk���Ub��V�?7�����v�/ƙ�=?���w�	�� �e�#a�^&�7Spc�w�Ҳ�9^��	ds��,���=�׎��_j�����'�q2�����?M/�*'��[y|*6���u��X����|C���F�G�E��Kz3F�����A�4}�:qXR=�ѧ�]+�kjKѱӦ�����J�uzI�ݖ����+ޙVC N@�=����nگ��	M\L�W��(G����k���U�h߸�L�>G�4q����������|_�ʦ�g���R�)R���g��l�\Kjd�+k*��69
y�G���Aėߧ'E�( '���4?m���94�U藚���wx���>�����Q�!� ��Te�4GӨ|�����a�i�ޒ�XD^�:p�>LH�b�&6�d�+'�q -D��Mv6#�K�������NrE�u�6ӽ
�i��c������i
ܦM��5�n��u8hI9��\@z?�2�bW�Q�\��K�ʊ������Qc��"檃u{�}h��	���[܉8{D�|y~�D�ju�o���"�5̟E+�!���!:���K�|l�7�o��f�`���h*?߸��	�
�#����+(D�:6�e��)�ƒ³
c�����J����"Ú�6�+��nbJ��f���}qצ/��D�Ģ�\!3~���s�N�F�f��7�\�)]�~RwK��O��T_
���>_���_���2�ڕ4��g�;�J䃻g����I#����j�o�#�\������e��ǌ[3��.���o{U4�y_�P�\Mr���?yF�:�/�5�<%��>ݓ0��{�igCF���1�V/���� c��Bt�G�i�UQ,�7���n< ������R~:N7��b�%�꣒8�>I�q�2&���V8�[�Y��h��ɯ�N�ӵδ\�R��l���i���͙�f$Z%<��M�f0uGpU_�w�8��ʨ�[�� P�U8j�`�Ick��YI���i������c^q�V����a�\�Ҏs1��56t8��SscJ�,����U���)����jw�>b������]Ee�-c�X!"w򲕶��xR���PY𥋷`�*ٷ�W��i]J�)o��	$�)o,���G�ՠd����tv{��E���=��@+$ب��1��lq�h#A<5�W�P@K���ރ���\�@Ȭ�6�4 ̸�8ԯ
QG~�����`=���'@�x�T%���ዝ?�Ƃ<fWn��3M��+m��S^�*�����ȁ�A�b���)H ��+'���Og)��(�-�w�"B���R�S�7��qYrO��w�l?�ե}��/�J2��c5�儵3O���7~,u%I�`�X�߬Bh��sJ?t��UE�D��"�<d�}\H�TL�	�����N.=��=�э���[]�؏ �i��@K�$��"C��"\^�5�<� (O
8;KJStd�6�sˊ1qH���l6�;	-�h���o����yʹ/&�~��ԍ��J%�;�����Ŏ�I[��$B�90�+O�4�+��~W�� �O)!��q���M�N�oX�

����ǡڿ�M5��{%R�

sk+1��?0��Jӷ�Ir����2g�cXug�w�����m�U����d:^�A�j<����<�;�N��11m���O��&��9=�}������e����p�HQ�x#����~� �G��'%��	�࠯�M3��'���	�Q)ج5��x꾧���+�P×g�IZl��� ����A�9�����{�#N�s�2�T�<�Zl#&#C���j�#��v0���g��R�f��[Tl�U�H?�Q�vr]-��2�YN��v��fQ�1X2��xh���*��]�C�չ��iP��4Y~7ar��@	P�6����4��uy桺���ş"����+�y�&������||pL���6
�{3�)�y���~��+�>@�[ ��&'N�I���"��Ư�w�S��i_geU���h_Vp6 ��QWCr���Ӓy�/��#|*ٞ�O��m�{<?���J[���uU�ބ�NR@M���1�F޻�l��#4~1h���[D*�Ϛ��R5���Sd5=?�IUw��u�"��\�h��+y��C��|E�پ�
�BB˴x=��th;�;��h�v�i��B^�j���� c�H�'��&�~�1C��o]H��ss(Mcp-���$��٠%��[dA�|+��[u��FGh�}$�S�Kjd{{pE\���U��y�Rē5ԇn8[�����p�$��
!od# �o�q%ś�至��Q��[�>���*�$�U)O,�*3�959H�?�4�a����9����MgM���Tjʞ�ޤަ�(r��[�ҫ���xg���`�q�ޖ�ZLHW%��ed�I34 WIS=�Z}ɀ����M2�6a7�f��Z���TC�0�w|ZE������R (Q����uý�@_5�r3o(ks��D~j�xr]�{4-s��N`�f0�Z��Q��W���@�v[xT�k{���d����Ή'ƌ#'�}��
���6X&z��ޝ��z�����
�y�
�U���3v��9eσ���ox��𶋄;/i��Ey��p!"􉕴Cg]9h��xh����E�ְ���Q�&���p0��S�MIc�y����Ze���qb�������*�i��u���(�p�L�����[{�Q߷(;�Ini�FE+Qpsaزm�ҷL��y��sݲmV��O�uq��<��`�>��'�K�E�,�1{�ȯ����z���mm�|�C�y���ɯk��o��䷬xRu�b��k�(&SyA��Ȏ��9wFZN����}B�0��0�a���0Z���؟=�ɽ��o��HŌ�*h�\�'�d�U�%~u�n�Ho0)�u�_b�{y�y�	3�0���Ą��y��G"�W��4��l��bY�AJ�j�� �y���q��<�)�y��b�����Ә�,��9��s�^X�f�h�f��v��EJ�%���a(�Y�Q�-��7�3s��R��y�)Q�%�&d�e���;0l��(I?���Oe5���;K��$�6���q��*W�M�ϫ���:-�q�J�y~�M�*L9�-�+�
��e�/M�c�QV�׀p̑K�i�Ǩ=�T�3F	h� :a?��)L�Ő<��fk�k���ڪ�ɿ7K,�7�r
{�i՗��.������e��nc��tl��S��K"R��t�6����w��K�`��Ո�.1��Ni���Q����|OK��i�����>���@���������Z݋�"�A7��J����?4�fr΢@�reM�������K�w- �A,9����f��H�e���!O�5��^=���u��_3����9d��z��Iɽ��E���R�1H>�'2"�~�'?��3f\�ށ��a�c�£�#�=&�G˳9��L��S�9��њ[j�TϢ+5�,	�f��u��I�i#6��^�P���
@���S�Q�4۩��nҽ��u����kDҰEJ�r(�T�]����O�|O8ψѼ�t�$zG�<�%�~o��N��a;�1e��|v��/>D��Hbs�vNZ(�0~�W�q<�S��5�uc@9�g�/���{OY��y�T�H��k����|Ȅ�/:Y��b��⡌8L�ӛa6�����1pd����q�$�B���'����Jp2"��K�~ �k�I^ʐ~��| e f�����v��XQ�1�����|�~�;}gȣ:���oW� i&�u�	�Ŏb����n1�H1aɣq�T|FԱ����t��⊧yߐ_4|��Ɂ��[����*Q} E�ݿnkY-G�+K|]*䟆����%�O�Gz�M3�,�W�e�`�s�}�.�[�]|鬘���ȧ$ 8�N�m@�O�g��_�\h�P��l�K,l��i5��*�����m�'�#�f/�T�I�} ?�w�V-j6�,�����C�dbG#�M���4� q�g>]@���ǧ,�|�~�/���VK��z�9�n�kЉ��c��^	��Vb;�����K���ڔ��$2K��v������eu-G�5X�*������o;��e�tx�Ο��� G ��zv�B�9A6٬�Q ^j;�ڛ?��D������	)�0��4:vw/|	�Rd�@��}Y �(<l��ڰE�ٗPc�xT�[Z6���k�q��%�(®�66�N.8�R�V|����m\��Ͼ�3!-(xg���*GͲnm\����t� ���ۨ�;ܗ])3Ӽ��`:dbT\��2��0��ԿgyP�l�� ���>�ߍ����J����GS��ȵ��=��(��g����RC㱉O�_iZ�ɔğf�xH��W��m���K��9=3!h�ɜ�{���]��֙x�<+�OUpw(����v\�s&wգ���PD���v#��S>��7*A��	js&�+�(��8q+ !,�K�J˨l�=�;k��y����F��j��^��� bb��"���T�qm;�=���<�ip�Mr�QsVI)/�;^��%L��5��E294jC7ܭ��CLx�.������1��?)��d#��τ	�t�Z)3�樃Q-6 <�/be��8[R�J {t�O�8m�D�P��~k?/I�o��^����[}��l���5�����E�N���7���ȒQ=��TG��"�<@�=�BW���k����������a��4�:��Srba��d�D�?q�V���~��o &��7�k�w�b[-��,۫t��D��	�7�����D�I˾��eeG�Y9x��p;�6sy���h���7��R�~�.3<�oO9Á.НO��?���9 �߯���T��p�R��>:��.��>����Md�j���[7)ڹ���	�l����?���)��$�3�R��S0����HY�$t����d�+4zC��?tY�t&nj~�5�tK��[�a0�S�|���Q��R���2r��
\ɹz�6���=4rȊ�E[Aլ������W%��R��ϙi�cYo��J7�|���⃂H>�3t��p��[b�*nY��j�����I3-P�����r�����"_z<���?X& }�._����������\�3��3���$�١��R<b�2����Q@�j[�If�zYF����p"J�т*	gH����,+�����%�4�R&6�$�-�K���pPɊ\������x�.v/�:l��sP7Z�M_�p��6�[F(Dg�g�5^���Lm6֘)9�%�e�Q����9�&���v�$�d 㽂ǨH ]��dQg�Ǚa5��(���ݘ��8@���bɪ>~�_Ih�B��"�AYK'��1�$�Ʈr`;_lˊ�r��Gi��_[s|���.��塤E~��D���e�~yqX �~l�F�.��?l�%�!�d}������r������0�p��폼�y��r�;�.e)��"p(.���?��mM����D0������^UZ���x��w`_��~��و���;<�����f%����1���z��x�&:
}g��6��[�.�ʗ N�]�����"�tF�i#m�3r#1�U���b�C�v��%x@�^�?��"�Q����Tmi��ͭ�
�z�_���~�}Ux�]�+
5ζIG'��T�L���6���ê���L\H0�[�g�7_<�gdq�Ԍ�mo���N�% ���M�h\��O���j;���u��]^j�	��[?��n�6M`)�턀pA*��<��o��BfsB�iY�Ä���8\PhJ��#@Y��D2P
���]�u���!!+>'�e
2�oW�^�Q�vϨ*�{�2gX��t�U�zο��V:��ykx�;LI\��hO�����Dsj�^��m����
��{��]H��羅�O���:�!��d�L�V�!:�+!7���wIH��'�de(�g�H}ͣ�ԕ]�����c8覴r(�ǜ��ʣ���轋�.�e����Ra�kF��P�kz8��qv�
K.�ǖF��E�iMZ\H�!�"rս��T :��ˎ.����	�?�	LN%�RWž����7P'^�(8.�HҸW)��@���C�zlW������0Ϩ�9�bH��i���f�F�i�7�38��	@���~�mB�KGR�@Ohς<ނ���.gb�S���Y��޽�K_�lδ,������p=x�٩wI�7��Z'�k�]�����;>��w�zk�$ ��Z��7��H��Ɉz�פ��Ԛ(a�!dPɋGIIDz	�����֐��J���F�b��O��/3���I�a��z���e���B7�79�/\u����E����\���ƺ�z�;���ʐ����-�YrF%�=�AZ�	13��冀m-��wo���a.k�0x������fE�4TH�����v�l�j{��ثcRg�'\����Y��}~|��њ"%�zʑ�,�y��k$�o��?1yv*�|ʄ�f���3�u�lǽ�j:Hl��}��@��5�c��K��T�W�82 � X����C���8��������N8�|#V�\T�]0���h;O͍�^GpN[��O��*������)�Bu��t6���i�/�Ay�l `	�$;~������\�}��K���*�]��R�8H�!����z���
<�?���
"��� �q���Tk����gks�kr)g�й��`��Q�G{c�J�}�4L�����(�Ym���'pTc�_��B>��_uY7�\�A��a$~��	��EP'��!e!�7vi]ڶ(V���@�n2���<Ѡ�r��w��7Or�p᪎��nS����WGTZ�af�8�lc�.���&����E��s��X������d�+�a��Fy�G��#]�ɖ�ĉi����*{�q,G;�{�U�ʱo�I�WC��Y���M#��ߴ���j��e�][2���?�᥆���'A�{�{��;i��mA;�I�%��/0t�'l�aW�x��r��*}��~�Y��V�Ùw%Q#[� �H����3,a���"ʼ`�Xo�������O����Dg���P��,Y�:�r]d���-��*���r��-�(�,����k#)������Ξ�q�-��TQ*kmZx_�Mzྰ��/��D �B����t���Ԁ�UNrbO�웰�Қ�{F�oQ�{��=���,�]�#{:3�[C�����2���'c���X�J��q����V,��Sp�kC��7����5�$�G���yeȂDsʪ�wFi�4r�׷*h,�JZ�ZY�k����"�C�0������"�&���Y����(v��RҚ��A�B�21Q���6�H��:�A�wF4��]R��]���6���@9���Ԁ�G�OC�v�O.>*�F�9���H��^��>�5:oFbl��Q�~� rTf� E���)ձ��3e�w��^k�P�-n�GIp֩�pe�{�����5��adD11�����,�=� �!��5�Դq�.t��F����m�κqh��T��<cs�2���{��P�!�񚵿�m�N��_���܁��y�S(�|��g���[ y;M����:�QƝ��|���x�"bP�03/%j��vZ'k�@9R	KD�����!/ߘ��m�/��-
���� q�r��Q��U�i�fD� KC˂�B��"� ���-���4�x9����8����ǰ7�aP�Օ������Ր�ndɠ�L��5=����H�nJ�u$hzL�|��%����@���yhnG�]�1 �%���R׎5a;)d�[O�!9�Z���v�j�7�e�|4霴��O�+�v��ۨg�2l�=Ԩ���t��7�8B .��iʾf��ya��i�o3��T�ܡm����:4��$}��m�_ Z����ƝN���4-E"����y���:!JD��E������S�������K�G;��d�,���6�	���B�x��L�Fʻ>���E�')�W9�ۏ*1�ڔZ�A�N�����b�n�B�b7�^��}�&nw�f����\;��&�le�U�d�����&���{>���VH2�_����y�nJ���\5v�2�̈́nH�ҧ�A�'�����|�ъ��s�U%�Q������/,ل�$�?�f}U-C�y�C�"�^H&� �^q�t��f��[���_�aF&�g�t�v�^I)� ha�OLY^�|���nKq]q�=R�'�]��jZJ�	�Fܥ�GY8ʷ��K���iбԊ�U��L�Z��j����^*��I$�$M�-� E;�������qz���V��:�0���88�� ��ӒH'�I��Pv�w����7�( ��${��m%���$t����K5�Oq� &h=��� ��CB���0�򌞼i~���.���~"�����ǀ�|�"!X���Z]�-��f�o����Ԁ���I7��ï+��ϯ_�m�B/����]�F�-����ݩ�3�h���)�O2�۰���j���Vo��VUk�J�,se�%�+�5ڥ��\Y��lU(Qy���m�����Oj�a���! baC�}��e�S7	�	���f���; ��p�)kIn�D��u��L��=��@E�����>� -+>ᷩn`�IX
..\W�˴���jNe-S���r�f=�
-<�ڵ+Y�{On�k+��X��� ��[!��4i{��m��`x]9e��%�N���V � ����Ep�/��E����'�H��i 4��C5���İ��b��jV��0���}�潠2��x�?��������5y"�1������U��M���Nv �+G05q[�����7LA�ŰK@���#��Zr�i-b��޿]BM�R����l#�`�v�	E1�+)W.��j�(�C�6�o�ْ`�T`�Z�O� FӌN���k7ݙ�*2Ф�Z-I�/�߳1���vT�P��ڢ�Q"��d]nv�_�)�0���ݺK�i1�{���C���F"��S�����F;���@S��ѐ^�>�a'�+}
*������;8�.���%�q�B�V�AJ=�?!ںs0���Df\`���$;�XP�c��K�Y�;=��ج�euj�5�Έ��4�xr�ߑ�{s�"@�`׹1�l�LuF�^yO/�U�A$�$�z4�i�7đ���q7�ۋ$��n+[kW��Tx'�xz����a�ؿ�_��.w�&	2�n�W7�&NϟJ�c��������1���OV\'.�hy��"�5�?vW���&z�@�@�
}Z�O��S]N�\�V��?��g{ K)��![b�E�1�/�бi��1��O^r����=��Y�����Ԫ�t�nE�N��B��˯U���s `Y��c]IK/��A�sk�FjB��죻>@�p�(h+�?�|J1�T��$4)O�K�|�F�D@�L���H�⮙ =�qX	f��K<�	YͿ���y_��0mBG]���zuQ�sՈ^�:y)�e>��I��]���d��R��4�<�M�PnQ�k�g6+*-G0JЀa[e[Y�A�!��`K����o\�I�����I�C.Ah.x��~�q9����݈�'�Y([��oW�j�#H�u�Og�{&�g[�ı5C���W@EE
�뜷E��G^!�A�M�.�#�6�T����U�V�b�
���$�
���|b���Ǒ:���e��$
|iJvVr�?�T�O>���d\�j��~����u������H�ES�g��n�A����BP�:�v��sr�R�$��
*�w���j��O1�/�f|}�8�	kxi/
5C��X�;J�p��ܢ�.�={~*�Y�4M�7��%%�{��ԅ��*�#7�����%]#v�SV�R����O2k7��sf=�i�pX�ʕ�Z���2C�,��U�ݴ�j�:���P�_b�n���0%��Ǡ�qiB�n���'�6"�|��$- ����S݈!HH���s�$��D:�=�y��!cpx�_ͣ�r��~��^_,�������B���Mc�F�c�BYK�:�ꅮ4�4�3�V��a}��R*]S�����=%��sߝ��#�VK't>3�#�y��i�d7"��h��v��غg�t��d�H3�7�	}�wno����C���;��ߤ[�H㜮��̹��`�1��d��$m:8q���=�cP��hLQ���}���Mg�@Ȉ騡ۡZ 
��0�Yǜ�sN<w�M�IW� �&%6���$�4i�GlG�@�K�څ!��o��{�|J`��M����0X_���R�������'�r~��/������ݝ�(�]!#�i�|SH7]�������r:���.G�2�C+�m43�9�i��Z�3������y��䴒�[~]�g������W�92��O�m�R�U�*	;{�Y,��G���L%�\D��H+�ׇA"My'���cC���RخRg����p@��Ł�mEM�! �k���e�w	��E���R�����Q"+�M��@����1�Z���xo_���[��A�2I�1oc%6�I��tna.#����P����Y�,��ds�D?��0<�\�E]�����Is�$��:��o�aB�b+18����i�]L9ִ�
iL��w&{3��2��8���)�A��	�����*��ƕ���H/�vt9i0BQ���,�D��/�$��$�F
eɾZz�T�M�I(��,D.�SW3�ob~���;���r4��t�����>Z�,Z�K��o�j~��Vd�<b5��¥+��u��v��/�py�����_8 �_�s���
����t`��y��5�&9Er�8%�������&Y����(75�=��	�a�*߂$��>1���X�s1��>���ʲ�А�%iIG�;��eQ����>�� ��C_���6�*�=�c��8m�v����rM<|����gmi��Q��?���c7�] �����rRC�Fj��Xھ
�	�ߪh�%+�8��T��hZG�w�θ�cu������C��� �G1�২:H{��UTyJUB\.Ɋ$�;�=���aH9�
1��#�Di
��a�L��3��:��hd�a����ŗ��=�_sKiʠI��JL%Iw�,�<'ח�����bRp�.��[?#��E~��q'���0 ��J��y����F`O�1�Q����%B���|��@CP��e��u\ۖ�8.em�{�S>�@My�b��զb:4w��x�1��8���-׽�k�Lj��z#����7�HC"�U?���m�3�V��ҕɑ��E�ʨ�8��=���e�`��h�$t(�Yj�#���du��K�T8���G�Ƨ��n�5���w�]�̀薝7���vg����1WTK�/f$�/ ������J�.�_r��j^M�X�Q!���"��G# HPBʷ��
L�K�b�e�_�F������i\�G}r(D��N���g�j�O��IH�=��a�{�i<� �z2�4�*��[���%�G�yq����E��! &�[\�k���k�3��V-`|c�� ��A����Wr5���e$���k�	=v��3R��6������stUS�_3[�nM� W���K��=d۴� ��m��5��<B��t`�)p6��F%�<}��V���Vh��<uv�#**cG��yuO-ؓٸ'� nu4�f�1�ӱg��-�	���溲�Yl�����Hl)�T��*����{z�]LK�M`��-l��b��{k�rꡫ��!x�$a~%e��D�:&�'y?�g�f)��N�т��x(�`�P+F��#mL��fy��y��o���C��T��]��X-"��|+�zc	�X\�y ��|�ka	gg��$��N>�:��ޯA�-,4�?;Ŏ�X���"��~l����Ys��L���ۖ�`\E�F����I
�a�sݞ���ԓ���mdp�mK\[�t���l7�����Z�����}ΑE�Y3u�J]��'j`�D��_4-JtQ� Â\� ���`s0�w�%~\��XK�3�@�y�(`�B�A:4�l���68�n��ga�k��&����#M��N�p\�7�?[��v����9רڮU�%y���j�#*���� ﬍ә�ƕ�8�ƭ�q���Qɐ���?�˖֫$(9>8����i����jٹ�L�^<c��ۺ���;Ĥ��bх��s˜'���$�� �T-ⱅÆ�bYIX��i١e����]ڂ)����*F���A�#z��n��ZMz~�5�IMK@���.�����q[�ʤ�I���7�g3a-�x���i�(��>�TW��������:���f@��T����MmK����4��L�d�1I��s_���.�����3Y�?2?+~�
���5�
kZ��A`��T��y��ǾD���sCLBd�8�܎/�^�g�*j�:���
��պ^"�/�5����0��c�����S҈!�jW��K���1��?��*P" ��C�<�Wh�N)[�ww�I����U����y̼�ߍ'*T���}��N_���C�0��N/í�@�lT��b0h�ma.�ۡ,yO�|��?��|���wOV���B�g�O�6?�cm5b����aD��9����'��P6������''|��6S����ΦZ���<��߮!�ݠ_a�0�c�-`�d4��@K�J�$
t�&x�?�؂[�ԙ"��[�oS�UQ��=�W
�����\8Y`HꬢC����O������7_��7�1X����gRBw����ͫ�*���9P�?7����n��c��LD�V����ۨ��i�\��4��qT��Q����VI��^��ڰ�%n�,铓/�5{g�b���/7gհ:�[�����"�֬VE��|E:<ϧ��0	C(y�)�	ߴZۏj� ���M���h?��+b�uL�ݭ�X� ��;��dÃ1�>!��n�:�\Y��t�:j���N������u�z�����o[Ҩ��j�f�Ș��jrc�P!-0�!��n�4U1��nɄ��聛?!��zVf� �@�x@Rޖ���X�a���M;�cJ=�]4����pn�)��k���-vť�.�*��M��DZ{�PRr;-��-4�0 ��9�WĐ�'�c�1���l}�8A�G`k��	�Y�Y��ōY���;�XC<h��~��w�_c�{�ϥh;��X:��O��b��V�"�r���� �^�/_ls�PP�*<�M������i_�Gm�F �x�lY�F�xT�ߺnv�%�ڷ/p�n����<;�ӥ1l�(�\��s*)fUm�*,�Ǳ��"n>���%����w��pZ����fn`��O�`��pǾ�'a15f�k?%��0��7����VeF�C��s+���'J�#!�h��ԁ�J �ƪ�(�C�[��x�&׏�!PfE���~�6_��k�2d�@HH)��%h%ɲD�$�|i�"�׷J'�ʷ����V*���� qX)���{�N+�&Юi�Q/I���%'-���W����rM��zUL��5���5H����{V�TO#�\��Lm�����a�ӕ�B�r�j�=����K�9�|��}��,�Y�w�	�S2�=Ҕ�X8�Pw�Ť�'f�D�^j��+&�KhL���( H\�֗�#��;�!�������>>H~�"��Y��}D1���#�l�S��|�\���E\��4#V|�ǦF����P���aZ��|"-[�VN��Z.�k�=F��&�FL��M.�&W�b%)�͠5�<Ɖ��ERs0L�W�s�PǨ	ʻ_~v��� ���'Lu��j���Mrhu�!���^P��ͦKdߩ�F�h��������rw�՘�Q����L�Yc;ƈ����?��j¡��;�F]���ʜ�����ՌL���y>�~��~���+i������,O^:�l�L�}3Z`�8�Ax�N�v.������ǉ�	�T`�έ�"����>�I`n�{-lFe�>t��vyn���4�����"��E%T���ƃC�t�3ox�ԉ���k�2ȳ���������`'"��G�j��t�n�.�!�Wm
���!���*��hq�l��.f�^M��,��u܄4D�^�p�@x,���J�H���}�m`pa���X5�M)L0|��c��/3�n�Vx�f Q��v�'��cu��A����o3N�#�6����&_���e�>U�`�H�~�l#�]�ŭy�chݤ��� u5K�K֌V�na:�k>�s�	1��S3����Lf�.�1P��)J��<�|�CC�&�����`ņ���*Cy�P$HfE����r�rX����N��2 Y,
��w��Y	��]�v�6�����p�����(}۝�鄉�Vlf����|] �ۻ��'�:�l>  V�p�|!���į��>gagS<`)i��k�7��y�	�	�5��6^���#3�j�	r�H��0&M[�Կ��/OT�ln�A�'1�3מ������w���� ��c�ؚ�
�8~:v=��>�z�m��`�$�����M08�m�詆� IN�����Ar3>�'e�B&k��#���ԭ����#tST�7�2(�]��g4���-ki\�j͈� ����&��}�]'�r܊-�$-�qnu�Z�}�����0��m�SN���y�28����_���#ҷc�P}췫I�kɤ!ǚ�(1�Ti����J7b���y_���_Y�[ ��&G���ޯ%fk��G�n�=��hD��gO�e�-����HX��0@~KK�22]�X�܂�#-�?�m�����r� �cDۜ Sa���Ծ���%T��f%ZW���敭��p�03/U���j�g��l鰮��[�$�#*M���y��Z�GS�ۼ��Ҫ�:���{��a��\�틼`��I|�ӕ`������s���<�""�/~�>�y�[E�~��n(G�)�yv�	zj�s�#�"��`��s���6*���@��v�n������c��^ɻ�Ծ�,�a~nx�_���3�DY�ʴ�w��hQ��ZW����l�~���O�R7	� u���F:�@��/��a�L�&�o��苙CGb��*���+7���rJ�=u�k%sM!�ʞ�K�*����y �wt*�۲x�j<�Zi���OP0��ɷ�(ʻ�vs��pz�(�����{�iy��9�.~���0�c�� $D���m%5s�$���.qPB�����M�a�>��n������n��ئ7/�͕i���WKϫ�M��U��߮h�ḟ�>@��W�yZm��J��� ��� �U�>X8����rk�s���;I�8^;Z�ދ��9MU���� p���uR}���u!�(�rt����b�A=m7�os��P$�����L�k{�~ Di!<j���<PZn��D�Ks{J���Slk�^>�ڮ�	�WN�}d�իͤ�\yj��0�4j8c�	.((4���k�˦� 9q�Nx�6��&7�oʶU[�*�c�"��Lk���Nċ<�T�29���r
#C7B��r�%�J2�qt*T�K���R��xT�AS�[9w�M�w[]���@���ԅi�pʖ��``��������@~EIQ�ڹ����G�OX�q#tҞB~4�e"wDc{�G�r	��N��]��J���Fə�V3@{~�pcѠM��e��>\!�ZV�%+�0he�}��?�{�*��k^�D�,0)�D�.y
��fa��Jw��gv*U-L�ɝ�`n^��]Zȋ���֝���[�׆h�;�[�Nݣ�}l��f�
K�hI�N R�v�7�`�#�_�~{���^b?~�Y�]ś�p����g1�H�RFs���@��?�J��[.]��@��%�b�q ��8�4@�U���a��P	�pkD�~ܒc�W].h9���\��π�wc���
c2���E�y���R<�Z�����QE�u���������DU�I���#�q2�>ƿ�F���<o���7�!�Ӟg��y�)�r�b,�:���d����PB9�TI}Aj�>��=�/���	��o� '�|��~��T��d9��T����~�݃��}��B� z���:!#����/m������Ԡe|�����}�Q���
E�8���C T1��xi\�v;r����݃�C��T6� ���A(�G#�{��a�mW@\�J-��p�Ҩ)�g�Sz��,0{�]D�*y������s�syj��S^W����0ԟ� j
>�����6�Yt�3�g 3��ع_�+���p��hM�f��!�=�`j:��C0�5D[���"�F��OŋXuߪB� ���HuԒ���`���X9�Hٕ=�%�+ԅ��Ò�fI�<�L{�3��1�[K
��%y"K��w�9�R�7��Wജ���x�\{�ۚ���]�i��Yz'�	pK�	������'��:��R�I��7����.i�u��R#-���-�E��&�!ޓM����"gC�dYl¢y�9�~�ZJ�{P�;��i�~v�&f9}��1M� an8r�j%Er��x����	G,R��~���[�/������,W�udV?3 (.���[+����:\?���m�:(���{h>����t!k���ZŌ7{-�ۥ��2����r2���R���/����:&��;v�U,8��|T�����+�XaL #��G�����=a���P8�0�'���:ur'��|��W�����7����Z�2Q����{����!�p9TW�U�֓�.Tb<yaTDkT��DD�УcF������F�J?KK�fky����[�W��2���Q4���{���:s���a���}�4�y:NK[)�n���9��h��� 5���U�����ٳ�(�o�����N���ׅl��8X�:��z��6Vs���$l���[���X��W�pq�Lا��1mfSx;REG�͸|��H�ͧ�6�u�Ҏ����oD�n�2��!��i�D0�]na�����M���� ��*�|���ǩy�|_k�n6��aI4�9�#�@a$'����&uT,-�`�d�-@G���l�y!�:9��0��}(�6(��Յ����/�
LW���L��r�G���#`���
���}!�4>�C �}`�����[t��w�7�솟�����'��z�i?����ϳ�1N����+M�P��~�q72�
M�S��`���>3��~H�چ�S(|>��kVs���`;�^�Qe��q�R߮�'�J��C0#S��8��Ut�l��_sz�9S)�ѢK>e:����Ur���V-:#���oH�<�x����!��e��Y��=�+�
@�o�#0 ��J� �^�h4 6�ͩ�%}NtO� ���ϩNe�@K�3��7g+�'$6]SZǌWbb)Y4�?�Ή>���?��N�vV�)b<6-��ŕ;��]3�Q���?�ͥe��q��u7��#(�L��!7�#�� 2���r���I�.�?���a>�0��`<�ٺg�
��KBކ��<h�Yn}��wd�X�o��J`�͕��xf~�|������aEܪ�ʸJ)�)� �qe�&�����ӆ%7R#J�'�}�� ��~r���-63�6�ç�c�hw�� �d�>4s	�B��#4d�P35�>����/v�?�Ym0�.��&)Z�f����'�W���lCz	�����rJ�N��� 5a��3�T���29u�qY�ړ����/�����j����?ē5;R,��d)��-|
��k�`Y q��dQ��g��=����r[9=z_�����fVO���NH���/�pqm��1 �Ȥ���Tb�p��K!��X�pPN\�!&Ӹ�
�'9mmnz�׏-tyR��x�H��C�h����ޖG~!�x�9�T�i�c&�ZV�c�>a>ƹ�ό���9�n����@��E�c�M�c���R�I���o��ܵ��V�'��Q<��'$Y��3u��~����0��n\v��}�U��Ԩ��8�����bad#��&�\xҷ5�ah+�=A*2S�3�*�`�b[+�1á3��z�R�(�D�4t�^��$̏Yx����z������ݠ�:Y�@&b�*�y!eȣbd�@үml%H@��0����QU���r���k�>@e�0�$̩F�>�@C���y<-�|-c�4 ��������'V���Y��5���f?&͕F��@m�#���C�l6��o;?��D�P\8 �m8!��b}���7sf��{>˹s�ϭ+ §dӢ�@f�d��:}Jd��z�V���1/회��.�������ۿ��h w$���ηU��S�!��|��]�ԡ=�Պ�H{�����;w(B���4A@=@nw���/��/\��-����>%�8?8���%FX˼����[�"K{�e���6�Ђ�E;�� ���Tݢ�{��S������~�w� x�n�=�a-��7|a��.`�`�bHbGCw[�#/N������-��s�O S��~3�&wʏZJc4�BP"�����!5�	���m��1%�-�a�K{V]���x?8G
Խ��*�&%�6�@���|����#0R�6��TŊ�,l_(������t�G,#/R����yjo�&젩ఞpZ.��B�.�A�?h�6K	��ag
*g(:z0�1��� I=v�c��{�Q2��F.���eq\I��$[l��H�P����<���m�M�'�ƥ|O��>�-Ѭ����*�}����sV�'�q#S�=�w�pc�䙠 �W�赦#�6�k!l�_��x��F4Fw���Q+	�Z?9n�44 �`�S��y�Kv@�7/!��m��&�����P�i�� �>�^oҀ�)�V���5Y\���E�^e'�O֜�'mmf󰒜�s�`F��+�}t��Qꞵ���FwMy���{�Q�>0�I�u:�'9��k�l��������'�<�qu���*%/;�Aۭa�l? �%��>�ċp�uz�x�Xg�-o��'u�!QH4�2��~���ٍ�򧁣��&=��E�l��� 0���יd�M�d]� 	��JOL����E��)�N��w�Om��hs��õ�^���>?Q~���9�I�Ef�N�_�t#\�:����(^	9�؏i#��";*Di���-��5��d��-A��"�����2�$���x�,g����ߏ�wh��\XR���{e���煵<k�����`OH���tX�C@��I�24��1�����k�6�l�u�b�i���I�,��
ڀ�C�t��aj�ؾ���.J}� �}��yΝ)�XU����BQ
�YO�Z
�WP-Q��1��q,�YNA]�q�����`��σ$��LPM=L0̴�5!�Tj�?����©A�ŇU���G�8*Z~;`����נٱ��opf�o���^o�e�İ���^�99��@M[z�RLNK>^���1耟�|��WJ�@�}�Ӹ���ӋG�Ad��_�a4�w��N43QC��x��	Y��Hs����\�sUξ�^����g��S�;��ˍ�Ւ.f8m�t�����_���"ڐ5Q�U�-�}�g
u��?si^"JĄ�'���q�lA��"z���}�nL��Ϲ�.�5e�Kv��}�d"U�)^h5 ��cIw�$U
�z2�oCr,Lmw�Teǒ��q��W�w�_t?/����+�u�Ӎytd��(-��oY�{��3Gx�`Q�?B� ��Ɏ��6܄�61b����~%�"�M���ٮ�~�ޣ��^��.^�Ǻ����<��qI~���߃$�]������3��	~���R_טe���D��V[��&��8Ƭ�f�/�.����D���l�o������|�8j{�w�,?�'����|3�j�n	�eE��.Ą얂�^m��61�������+���B��-�Z��ؠ���� hȂ��fSf��;Ǔ��ޱ�<a�:�k�X'� g��c�H���R� 1�7n�Q�Fp�R�$+�i�G�:�jB�=���D<I���:������3� �1L��	,�|/��3bN�i�I~�X|����#�
^�Њ�S|��]�pW��f��T��u3@�7-�(���7�L��!y��m8��1�+��I���T�mGUVM�V��Ϳ�"�90���>�����h�Ƥ�,@�{~�c��Ц��L�Z�����t�E��t���U|�����z":l���2���0`7#��Y3��2!t�@1N�.���������CH���/�v���4�/@�9�[S��%L;r3��;�2�l^|�~�)Q��T�ά�5��s�:K[�[�sN�q�mR`j3����/2�O3���O#Z���!��ۺ�y��"�i�ݞNRJ6����/��n)16H_�j�j�a�w	W;%{J��9�~�l��TYw�Kf��U�~�p�zB��f,t:M�P>���\�i��cWAt�@��9l�������%S�3:�qSu��l
5O�і+�?jA�kؗ��#9�g�赩�c��{�Ѽ�z��{��A<���비�%��m����P2�ËE[�Y!�\��q����y��?����[)��f��>Xc̖�F�.8_Z|��6W+�3U�9q�(��V�t��O���E�L�x�O���!����3���!%D�x��=�I��G�,: �����,��Z���gm��Ǒt��ql��R�+��"/��f�T旖_!��$Fwn%�^r��Ě#Ak��LhR��G'N�y���mW�'3}6�u2֔G��w�_r�7���N�cK�s���>V(-n#_�_��É�e��}-d��ףּ��+7�N;���qW�&R6P�g��P�����Nv���̏���O�U��0  ���KISn6��b�x��TgmBY�Oc~�������j.�
����_tvı�U�T48I�N(�AiO��ſ��Sv-���}� 6��6v��L�MYu��.��[#�����B��(�-��;E��"ʏ+�~����Lw�a� �`��[�<)�s��Ihy@3,\�;0��-\a�yM���SK�F����Mj�u;I0���QI�U��}�elh��vEVQ�Ap���5�l���S}��ᩂ�E~f:���)(�V�ur=Z�(�˘7�����Rt�7~|FpO��ɌÙ4�(k�Kc �!�� θ02�p�C�D_���)�����h���+1"flU7��������)�mB,Ov�~0�+�r�ߴem�̨C��p��Z}���VE �t`�-�P2��=��q�R�b�әn���	�YS���+��� z���n�K广��h��L�!��p�F�Cn1߿����M�~R��P��:ݱ\3�E�yUp��ͤ��.��I�S���\`dQ夗#�u(���&[P��_��x�t����nS��p��E|���h��3�����s[0��5�S�X�q��FI��?S�r~n5��w(�m��}6%�T<Z�:Y8zw�N%����e��4�
 D���\��z���[v��eb!���7�H�ѤP�6`���&��(L�K���y�c�/K� �.�)�/�؈�7�{7�ҡF����|��q>�,�P�Y9dX�1M��ZxW�
�h��K��XC�1�!��G-��o��eVaB׮#`��!�t���;ŲVh$���0�pP��ε�.'��U/��=��U �>�/��gi��+�I[�}�1������5�Ֆ�hq��ڶ<"J:���+[�X���6�|1�G-=��Y�/v6;ʋ{�!BO�ďSyC�
ti�K�(���]Y����p<�|kO��8�J��?]�1�]xZcF���GAE����++]>����L�&�����o���O 3���;���!���qP��"�L�>}*DJ������"GzAE�� [�b[SeYy�D �[�A��kr��5�m���d�&8Խ�.� �z���і7+�l,7�)u�B�W�*�=P��"*�eg|ޥ,�F�H��`ޖ��VKc�z���	U5���>��{J�	4���&�+v���]��}���I�ԿaS;���`��[ǃ�=^i�G���ܨx���
�l ���Q}�Sf,�n��1���D@�^��o��;���jv�ףn����Va�H����l=�
�����`4�;��3��f�YQD�~���d�hT|2_��k��W�˶�?*B))9y�u-9����5Ǎ��>�|8����ê1��0	J��N-:�ݶ�'�f����v%]g��w6��k�"�����X`n��Y��rē���X������%�8��A�0�3�%@T��ߡ	���򥇑��Ƌ��'�`7���r�����4�u���:8j�l�*nm�E�g�a5�_����;Ѽ��I��1�l+o�Z��I(�1�b�F���i�=��>LQ���a;���}��]��G�b�R�b��k��?�OTd���5����F��h��4Wor���}
�w��' F60�@�1�-F�HN� �2X�p�������;9�p��i,���5I��`+$������*4�\㒑2D;�s�1Ǐ����=���ٲ���i��x�f��8lX/��/�҆{ԇ��A	�k��Y~�G���1��i�j�$B����!�F��r�M8�֟�� u��!�c��Iϸ�jeD-0��v6�PA�U�����������������&.EYS�,/S�` 	�����-���Q>]X@�#����6M~����м|c�ZV$܋ƹO�֗��!ȏ0��rq�>y⢸���u��M�Q�����8ȹ
�se/�׹�b���R�e	�9��4\H=�d�o�G�dL�i�o�|�+ɾ*�q��'��
V�Pu��9�XnX�����)C�;B��S��ǯ�����iT�g��i��.�wY<�2̸��{8��
aNfӽ[���Ӻ���N4��|ǧ������]wND�x{��K R�P_�q�zye�fo���z��S�gɤ��S���-�|�J����+I��+%�+���⸊4�Üm�3�qg�%�Z�: =��K��~Vb����Tt�~��%7��@u��?�qח�|+������N����qC��B�^��C�C�j|�������b�
\
�#&�,��꒍����˽기jJ�O����U��9����O����4͍�q#��҅/p:5a��X5��7�Չn�qiy}>�T���K@�w���S�_m�gO��!ߣ8��3+��(�xd�l�"�>C����E�n�䪷�K̊�|�4U������
�<�6�@�ˑ���������)�����m9�F�xY��D2'��u>��.���d�' �].�ˉ&ܸ���T�R�|�3� /Z�����K7|=�q*6OZ��\R��p���&��y����k�`�٦M�z�g�ɴVy��<��&�l��
W��o'2��%Z� �˘�B�4̚�5��_.^��f�Mz���3N)��6.�i�-��1)T��i��!�p�M����G6Mb���n˃~Eh�fз��ّ���jR���Ѝ�h!���`6Z���[њl�������\Id���53v��H�7�,W�6S�B<��t�X����9ؚ�G`ڣ�&��T��z�>��ҍU�r�F�z���<~�u�!@��wj�){>\X%�Oa�^��Z)�7�a){K]��GBNh�+�*%�/��TĎ�����=9)N,�<#I9���I�oA;)��^ִ��� �ٿ�?���h�+��io7#��2���$�	M����ˣJr���бQA��5���+�YI��Y�~��Nh�|4ǡ݁�<�ő8C���|���[�Se�����z�r��o���w������@�:*`�@p=W#�|�����f���w2S�?�E�9�q[�+qu��ى�ڌ�#�LBf���P�d%�M����+�qw�z��9���Ⱥ�� _�x��0`�%S��w�m�3�9BwG��Wg�{tq�Ԫ�p��xP���I�5GV	Ϳ�.R�h�,ٴ��>V0ǆ(]/γ���K2t�.Hx<V�x��o�*�_���4֩m{U���~`�0��o�H��QD��8�Q��'��4�V�]HS�l��$����J6����i���i#��9A3���:�����6�B3{!��#B4�qS��&��6ceø^�	��O����>�ˆ�zfq���d��b�=�yT���<ό@l?��G���
�=�|L΁a��bP��R8�M�=���bc�"'8���bG���R{������ǔ����/����}�j��J�� ����� �:U����׋%����Dph
|�$v(���K�E�L����l�ÏT�����B+/��n�@q�}7�~ጹcϡ���Q��w�W�P.�)#�/Z_v��A<`���*b̷EN�a�|ONL�0o$�#�z���YS�VƼ�� ����X{"'c=H[���1}쮹H����*��h�0�L�D2n��L�_�h������ݩ}�%��E�#�9%�o���v1�eȾ�_mظ��9�Z�,��3��ً0#�U�{�TKL�ϖ�y2N�@��6�����o�j����"��s�{�o�q�e�hL�s�!���+P�z���hcK{����o���S���-,�kv�d�c� �}�l�9�|�#T��1�V�"۝䶉����W�q�ӏ�8���K��
��H8����3=������p��p\3n&�/���H���BW�W
 ��`��V6��^{3����Ŋ���a9$B�=0��~��g�Cf���P�g-�'���}�y�2��s������M���XV
�D�i�k���?�PէRu�����L�znZ�?0��k�`[��9���k7��ۉXKE��n0����;V� ���މ������wxk���}9-�6Ge��T���+v�w�ލY�1-��-����a�Y�N.��ǈ�����a"]���/�ة!h ��
��A�X���0,��'H�����m�[{e%M[.�`�@��.0��X��'4U���Κ�V����ؠ+6p��b�$G�� i��M�x(���}���ʩ��D�Шb�9]���.���`�fP������K��9s�Uc��"_]_C@ ���=&��������L���*��@�ʉ�g�p�tw��.�i��#�g��!u[I�wƩ��me.�E��+�'���Fp�ciO�QiK	�
��[݀2����)Idil6��S�q�X����{�.J�re������z8@9t^��@����:���#C���5+U��jL����qw���x�Y.TbJ>����h���:�Nd���|[��v����}�O�m8�-<a���Uz6 +G�o�[�N�.�* �϶:��ۢ^��[�껋_k�(	������m�M"��`s{�o��lek�#s4�SD�nM�bݔ��MAH��U�>{�#.��02���Hj��/p	��ӧ?҂r�\sr"^{�0�_�I*Jƛ���ٶ޾
K�ʸz�H��-��~Gح�d��G>K^u��_>�闍F�t��fɀ���{��L���lL��>�L���.���~{�J��@��J8����hoH��nC.�-��P�_o2@��Tb�ss��j'(�Gޗ
�,�&Ap�a�~�s����cR� � 9��P	��Sz���A-3Y�ᑛ�v%`�KMT��%r�%�t6�n�zZ�y�����|��6��^/3�׌�����'m���bzN�P�]�sJ���]�Qq��2���=g�9 �5��	դ;������1�4��P�@>b�^��I	���YL�������y��?qAJ�ji$��H�t$��P�.�d�������9Z�z,(%���!�Q;{��ڷX�ȑ>�F����)���ZN�s�iR㗳�v���u�"�ț���"��4�y%>Rӽ��<�!���F�T+ϯ�^|M��<lFQ��% �5�(�Ģ��;�������e��mB��t�~1w����wt�Q�B��:��:���N��t�p���؊���~S#�+Y�h`z�����=���]�r���t@a�-���3_G�ڪ�[��y�����;��Ֆ�V��JZ�fN�l��bz������Ʃ؇�V9�ʲ[���SK�>�?����Hӗ�2ɐ�*PdKEGw��W/@a�i�S�[xO��NԻ@�a��5�*g7RF?u�FvP��5����TAP\<�
�,:c���e�Z�*�b�R'#U���s舆ǎ��k},�ѕ����C�ˣ�S�y3���9�Ll��o��?���SI��6j �#>W^��`�#��v����MQ��8!Ks���#�@_�5�)iL�Q�}��O�������;E���y�,	�q7z�;j>5��!nZu
�	�=y7��P�3� �m>d�6�u;D�VU��#��F�M=}n*��gP�(	���q���x�%q#�����#l�{�_�犅P,�IX(bj��b4q�Fɧ�j��Z��Q���ay���m!�"��D76C	��?'o�#ô5;购��1�d�>3�ڏ�Ŵ{��ݘG7��C�������J\{/�VV��CM������1�M*��K/[�J{�մ�P)��s���K�4"*lfbkda;�V�Q(��9th�̂b`]�L��[]��>����������,P�ֹ��Öt�,�W��RJ��w�S�jx��c������9{��M}�KG'h���V����o����e��dV�!؜�C$;�����h���`����ؚ7���^H�����M�������Y�iCw��s��jR�7�p��C~�9���l����z�O�q�:l�({��x�Jfl�Bk�w�c~{:��б%��HO����[p���f'�W�[��Z ��"D:���9)|� �~)F�Cߙ�V��xCQ�<��B��z��Q���]T/��?3%	����A�q�x�D��)r��I�#V�|"���'�!���s���U�<��K�u���H���ߥ�7��'[�>mtţ��t���a��]�p[�&��ː��?�n���H|����w8D#oeh&��b�+��`S�
���85|a���&��+|��pm���O��i�A@7��Fb- 2�$�9
�l �O;;����p=-5����F?���n�����S��es2��rՄ�GM�o�q2�c� �EA�Q8��à_��В��g>�Ǝ�hL�B-ǩ���T묾���|��9��X�� �:�5�b����y͈�M�&豋��(�rOi;a�\��u���;-,9�ڠ��ee"�d���\��@MDG,���,5dN΁�Q�-[ƕ?�-��+���Mb� �oߺ��>_%I��q�N
�}�7��O-��M\�n���y1#4�\_��i�nXW=��x��M�Y|� ��HR��e6a���Wݸ��x��\�7���l�����f|+?�ƃ���5鈂���mҶ�1�>ܡ��7Z/)�cÞ�����?z�j���6��4�c{�OM��R�A>~V��4T�38����ٛ��g>X�@D�V�`��h8�[�y� �s��}���԰� �˛c�;�D�^����v)/Dk�_l�O���;h�3\ce�=:���C�:O7	�z�\��D8d�nI��������w���^=�T��`�@|�[�ʜ�6���䁴R07
.��@+^����t�@��5�b�Y�V4y���>�
����3�蟺Y���:u�-����M�ȁIՖ�DC�Z*{���Q{ַ��R	������@�G� �X�.$�ۓ0�&����.�ࠀU�q�lRk������A�iG*agQl7Ҧ�};��R��4-����S���g�H��i�ܰߐg����+���_�1�m�����P���E*�mM��v�3[,�� ׭�[���7f��}�I('�����*?f�=��r0�C��g��'��&�����Js�N$}��ɺ��Q���۬��<�o��@5��фѻ�'3N��3:*��X���X��:P��>P���'E�/'�Pf �c������.�����;̘�Dlc��"�i�X�:�i����tnLW�=�t�dlq�KS�L�Z)ޔQ��Z�(}ǣ����^
K�@�ם@YА9�sVe����@EM��t`���se�F|xHcx�/��4��x����֨O���y���<ZN��is9*=� � ������tx�1f`��6�������4@^����/�h�5�?�-����L�H�i�`!�Q���(eS�a��tZM��5��&�o���'_�qZ�R���Dcu�=]I��4AVqX�ZVSۿ[F���ӣ�6�����O9lP���"�u[P��(	\N�cb>�Fحg��l��A���v/L����L�>@��f�{������s���7cC8�����q�bw�/��l�f���m�,���:�܍̈ј��9P�x�"61.�Xd�y�]����a��P8���bۓ��q��㤤����};����W�~y$z&y�>D�ī�~8���ǎ-���uI���W/n����+�#J�܏� ��a)����nJ�����.]<�0Ƀ���%�x5�Kc�"�#$!�w�y�f`(sj)0����6��d��?�����d$��*��R=f.cG�{+�����ʊE�2{���)��� ���}/f-c�"6����:Ȅ����W(
~�mUU�5�Mޔ�������/���3Ͼ��48��W%����A�D�%�V/K�G ��`��,��;y]<�"`��(ݵ��8ߗ���������š���w;�irS�4��{d��u ��?���Lτ@��Z���<\��.*��ld��w�|�[R��k۱���s�"VWC�0~�L#�SO;T� ��A��W�E�������@�3�f1<+Q��6�,�����Vw_^*�z���"k�
�����pg	m�?�	���z]`dDoX4-�M5(��L�9�P"�v֫NT�M�g���&h�dʾ�	=2����6���H.�/j� �:��O��`�Y����=&Mm]�ηR'��m (iRB�;�qW�o�w}TTd�ZN>���[F�2�,r3�\p9R���t�Di��;����nK"Yr��@��K��l��T�,��"hG��'"j�.�0!�=bY&�p^�$�c�j�'��m�g�1�ZCu����:��ր�;)��X�lq0�G�!�*��%˨��̭H�L�t���'ᆞ蛙�#9�-��+�4�4=����oP��Ld�5Z�S��Q���D��H�ȇ����U��6��-�)G����#�b@3��"Bش����[0`n-��*9\����:�$PJ9��N����	c�xMiC��������T��W%X�C�ah
Iܬ>����	%��C��(+hݾ��(����2������]p#����0ZO���������mi�# ��]��N���`�0�)&V]�(ޭ��Y��1/�Q�z��F�9���3�`���VP{�����d9�PB2l0�dZc6��ڏ�?Zp]
��>t$G_���y�(T9}�U*���> |@O��(f��V?�6BhQ�(ķ;��|6L��O2d�&rj9!^t+ã��Cw�����PU��2K.���/=�Kˣ���7��	��/j��g-��2Bk���QMza�\�O��9�4 ޑHb�5�$��*K�WF~�����Y��	�#ʁNņ��/�k|*6G	�;��կ�m4��`�nB����0#�� ��5�8���f���chS͌�զ�lu5 �l��z�{�`+�m�a*����lp��>t&����S�E��i$��ՈbLT~�]Q�@T�\2�<?L�E��9�
Ar�u��� 芸,���@a��8��բx��d������<Ȝ���讉ȶDQz��3������94��!��	l��=�%�5"��
��f���d�o���:π����P������ ��3�}]���N���K�]GE���c��|��e�3����mG���Mi�	�9�c�m���H`��f�d�.C=`n��4&��^t���5�(���b�dgorlSK��u�puX��, ��d�t��Dl�s���ѡ|���~�X�О�Aڒ����i}}�eݙ�>A�6�0e���_Wqؚ�z*^�1�"Y>�c�^�#٬��'T峭*���h�p�Y�+�J(��`	-��!���yV�I�$��%D�Iq�x��H x�obڱ
E�(�
ގ�&
�`G���{�ci�,L��T��u��Z"�'�u�0�N�a$�iD>5�$8U"���:�c�+���O���f��}�%g╕�)ͶJ#Ԑ���I���.�I.P�*/L�»Kn�����`_
G�-���Y�aX��K�U� �-�?P��3�_�C�t��}f����W�r*���a1@�-���[�ܨ2Kа���^��z�/��J����Zk1+W ?����S���쓊3>��_:��j
gu�$q�Y^���h�@�����'�W�<�mAoq+~�"����YT$�L�ͭMu��=@6fZ�j��I�o#�_5�l\HF$�����Cp�h��J�.��ҥ�š�J��`��L�|0]?<(�L��Mb+ņ��Ԕj�J��/j����A�Ǧ7. �ڵ�d��T�}����b�X ��0���-JoԱ!��W��#E�@�0!��Nr�Y��L�%8�
u�Ap�!		g|HfA�
H*Ӄ��T�������he�dW��]���#�A�J�Bj��;�����+���e���џ$A)CvQ$�3�#���u0��AJD��pHi�1��.�$���L#{�4L�{�GJ|�Z>�Ue�հ	�����&e���5�k��%�����7S�8�F��bc���~���f��"Y�\��[^M��+D��'��x7P@���)T(0����)V��޾h'�Kd	��w��^�AL��Ŵ���j*�T���Kp˿Ms������3��|(�89�[ ��Y0.|9�}��*̰c�wՄ%�S%3�WV���ps׬�i�Q���[��?�ٕ�;=�꿒�D�lKZm�fR	$.�l	]�'�)AU�#޳��_�@-�������cHd���M��iU�]��/��e��R��Wh�P?��Ћ���҄U���U���2�<F�*���Q6W�*�ֻ	αw�pD�У�c��a�'E`;�'�<�u@L����#���)b�7���v�u�5*{i�M���xv�*�p��Ͱ����!�zT������ױ�f�q?x�w��vRmҗ����=8O�o*5�{����]�U�,���@�~/P+3�孲D/�]�yULAm��E�����ZJ��$����?�?�&UB�
Fփj��$�d5�n���%1�W˻LMRl���`�v&�b�^A_m�}�Q�2��=h���)��l�,�j�ԙ�A=�\�Ak����k��̜��^�<"�m�\p�B�搌.� Hg�|PK:�J�?^�w����Q���s����Z���_(�e1���cP���X	&�C�L$�y�q�#���l���ؠ��F�	)��[ˉMOW�LjO�	g��J3���j����^�֑c��w��]^� 3��b��Wa�"{�N?��o��6��xKi� ]��,�d=TdוB@�k�ɪ�>��1%�@uǺc�_���+�n�V�i�qF
"(�3jz�*`Kg@{/_>���5���cx�i�f��X�m�آ*��^+T��$P/'���g�8���ӿ-�]�]����`�&}:0����z���}s�Į�q5{�7�;m�ՎB��N�a��.�Lja҇`qZ��Ry��X�C���7��bdB��jm�O�{�kYcϷ°� a�>[墸�kw�Mk"?i���"����Z^]H���>>]�J3_.n&��Y���m|�5B�f�67���$�;�8��H��+�@[<E1fp8��imE�n�J5\j���]3���W��\͜�bJ)���}gE���:���6wi�@��#�Y���2�<�i�q����q�x��+[���#6�t0,S�r�?i�����;�ϐ�<d�*�5�v29>��G�	up�	�����i�^��i�L������������DkjU6>A��0���_�{>z�F�4t��C�pH!Y+e!�Z�-l���;�5�w�uޗ{�!��]wSSD�3���2��������ìe6��Bشw*������\�3zs�߄#$����|g~8ۑ	2�Ra�BKÍ�+���q0c׺m���T4�.�HM"T���o��Ei M�q�ٺ���]5"�sɛ��^�_����<����8�Ni�c1�61�����8X�n��-1U�Ț�M]ļH@;�4�k��W��ä��e���ȏ�	3X�U�]� S���u�$�ѻ��q@�3g�ħ1;�P롫;}�I�I�����Q�џB�}
� �1ph��� //�����e�����I���,T�j�D�<������0�w������i /����S@����i
�w��۳��?��s�JZ�_?��y;
�p����}4՘�28�|��l��dEF��6���W`e�LfPKO��Tc޸����]"��*Y��\]�"ڈ5�+�$��x���уjA'��(`���އ�G�i�H�2��ڲU �)y1�k��b�I������[X��'$(ee�2�L� R[m=!�ψ^?��,�Ҵ��#�����D~����V������V�������1������T���L	Z���X���>S#pp��Ѧs�YWkՐ�eF���6��}�E\{���v��G�ojD����}�?�ܚ4ro������KK���
DbB���.�~w׾S�)1�v��D!��E��&��}t
f71���l�؊�I�B���הW��¹ͱ]و��zy����Z�?][�1�/�D���Hf�c��n��^mH^��U-�L?�������͚w	��X*�䄝i���s�M��A����@�U��$��Æ/�Su��<)
�o\R'[6tJ���N��I�xF1�����h�Y����dxeQ��@��[�/�I��$F���+4EF'����J=N���L�˯�t(J{t�vY0|�^qZ֍�D*� ugx`h�����U�ƙ�_��Ε"�8��2]�Zqϥ�`1O�M�@��XO���evQIh�v<�����j�9����F2������]fx鴭���'��\�'F�u-Ib�ޕ9��A�|�B�����4�bsG�s�ݒy�8t\~Q"~#����@����g�TaK�#D	Ն�D�?��˃{:�Fk�d��h�d_ �
)3CR`"�bd�-����{PVE��X��ȤMJuOmG����щ�z���P`?$�rk�EL��a=�VVl��[�M�h,(���i�g�a%�OH^
����I^��\�J-+ݪ���pb�_�MиN5�؄T�PK���\�f7������!� ,쁪n�'#���|.�ڝC���kW���!ʞ%�2�&q.��'�d���]�l�$�^����� ��S[%�?�n����0�:>x�����
jT���A���h�=FS�R�P���8��Q�Ԙ��nK�Fz �E�_X�,�����'M���?��$�Dr>G�ꃁ������?G��B���&6�h���+��p��'�`0�p;�ϻS0�Q"�m^�4�����5��|�B���џ�����՘z$mat��8�W�S�`Ԅ��������[�S�(ʂ�$zE&;��e1?��0= U�Up�	A��nq���v\��
�T��Ryn���'�g��1�u(%��*k�Q�����-X+��Z.�R�0��/��`���^h�sڇs�(Pq*q~	t�t�+��&��CU��Z��%/l�P�NN�}���>l�����IE�i��5���9�mn��%
V0Rt	"�'��|�Ap�L֣p5q�YM�M8ӝ�G~���Z�?^���eg�߬�����o�P���񶝄�I Ģ=����*MG�����L�5o��=�S��&]@��nD�l��t��@��ߤ�o�������g��R4&�S@[q�����a]��U���A��g��� v�}g�W��T�UpFM	� �3"��������8�&dƳY��rG(D����(ߞ�HҎ ��|W���B�	@-�,]���6io�Iܶ,�nP3�T؎�ı������ZdWu�G QZJ���X~D"	5Np�WfZ0"<d���S��Ɔ���S���PJ��^^��/1&��*�߫��1� �T5�tp���Y��M.�U�����*��i��7ȥ"/�WXh~)�[�B;Uk�NX&�,"Aq��?{��wXZؕ��B���~E� �>%����=;2����~�5���;fu>>�����	n��X���{����;�tKڙ�&���b>h(cۅoC%z��_K7�*.D� _�́�?l#��z<��̢.R�U�]��; �s���R����ZvM��&tp9!�����:�t*wdvQ���F�%J��ܮ��p�:�5h^�5�&e�5bxC�l�2I4'XϩA@,���f���P0Ƶ(�/��H�IO4�ڶ�PgohC���?^��@F�W���f\�F0p�s��� -�)�@L�)��Hc��4�WRM4�v@>([��g�8��y��6���?�P�<T��k���I�Y���0�Fj� I�]c��:'J�2=і�'��W�"�,���[�dn��s���(��r��J�+b�؎'V8&Ш=��G��Z�J��#i�wr��vd�5[�
���W��}i��z)�x���K�n<!fc�RO7a,�D{�>�Q�m���������l �UOR�&��Ç�#���:K�����\*':9���#�x�	� �։*����%3�X���f~."�a�M�Lzv���Vzذ�O^o�M2�ڼ��1���z�&dFF��Vs�6�^΁�r�Pp�B2`��b��bML�KB������Q�G��%�1�b�R�eO��#L��ۂ%N+���{�U|4���+I�&6�����"���dB�u.�"'Ov֨���r!��?�Q	�}�l�	B8!��jھ;9����q��Y�WM�=�x��D�R�?
.��I�RL%t�u|���"������m��߀L��>9���>x�9&���
�zE��"�N<�N�|�JJ)�Z��[�Z�9�5�H��mEoL�:a�t�f3z�8(V�~)���I7���[`N�Z���1�F����c\$�м^�s�W{��ۗ��y�0%���v4��E�rբ���{P�i/��`-a�?��_Dd���\>�*Fy)�3�w���R1�&�����@��%�Sj8��|�;�@�_��o2}㵜��\�q@R(�1��㗠�z���ĵ><��(��2��#R���������\�y�l��g
Q .>���Y4g�~��[����<��ߦ�g����Н�X��X��3Yb����9�FWj�URRI��h�(�_�Y�PL
xH����Ei��Q�GpΝ�i�U�H���! ZP��r��+ĺ�k���h#G�PF�F�ϡ4�q	��L|:S��=�H��C���q�<on�8E7f����%U�u����P4��
�z��K���W�Z�"|���(���yi��`0Af4J�Qi��\Ky���ޏ�Z�n50-E�!4Q �X����
(��7��f�h�x�i^����c�r����2g�EH��0���7���s���3M���Wy$T�Wd5\$�V�;�7=�2�ꥱ�}����Z�!∦��P�؈皠�� ;���YR�Xzd􋈎Y��VCJ���k1�ּ�������u�+��p�k��$4l)i�N��)��A�L@{���|7�������RXԍ�K�Ƀ谐hd��*�/�y+��9�ᰠ#Ą[�}�E�<�	{`��TwFe�h����}G��U�@5ۢLB�߬hwr6��3���*���h[��O$p��{d�������:@OgrgJ���{<M)\�G1��R��t���DL�Bu7��Z����<�5Q�CE��Q)�Y�bE�!����?99�dw�+~İG�j�
�r��X��ZwH)���4�/.��:���:�9la�@;Z_��Wb�+23ѫ킹(�/E V�m^|�ݑP7}�s�`R4ߴ} Ț�q�k�h �+��o������9�3ִo=q�ۏ���%p������ki�[]����ۡ�����g�~ z� �e�������ѠR�Q�[�v~��e�Ğ��1�=�g?�����W�-�v��?R�[�-������o�Ţ^�Ʀ�Ѳ\RՌ�:غ�5 ���u����YvY��C
���noW��L��OZ]h8�&��Ĝ0���x�ε����8$���Gv�:�@g������yS"M�u�m�?���F�k�!�/Q�h�l���M��-�$5��r�<��"�B(�P�H��
�bé7����=�E�0��5j�=$v%�,��Ļ�.��)��I�?���'TV�fa}�)(�o{�M�PW+����ܰ�6��&��c$�>�3L�XN���)���%��]]�	�v;�,���O�Fdq�dS��*�G��X��}\�����2�����=��KU�A|���0�%ڊ?6n�U�!(��[��I��K�Y���R�ȝY�|��Stk��iZ�`|��u�F?s�f�R��#�Y�?]�;�)P,A�-O� ��s��ة}��I�)Ue���t��
��
�:ny9�u����J�쇸�����xN���f�ߕN����@�����fH�h̙� �_D<���+&_�Fcec��� Y�N��r'D��5�=��l䓠o�љ�yH5@�n�&̅���S�d3	�>�
g:�^�i�	9'��96�Ә2�\["�9��r�޲��}�������J�v
� ��۠0�i{��?�6��+ؽ��"|V�-,� �Lk@Tt�6�U�a�͓Gt�l��c��&�7~��&���d�ru��W���qt�q?b@��t�|)�C�XE$��O�E��-0P|{f
@G��=��n;ߞ@e	��W�Aځ�l��"Nɤ=E���m��M4y?�2<�ln/N��S�J���yz��`�S��d(�3� �3�|�s�ˑbɾ�`k �d��.�lB��P.\�X^��M��bv������l�T!%���a�y�g�X(o>��%�o�n��NM�\>w�I_U�Ҝ}�q_����p��3�Ia1��u�G����� o�M�`%�?8��o� b��/��E&�}j��%�팸�O��I��!�gG�h�`�5�=�d\� �K�}�^aE5���P5���֫��Y�B׵k�H�w�����O߾'@�C�5�/@W�#们��E�3��U�E���&7�~�˃��t�-�I��#���3���)nR�u(8}Wϖx9w���!�v�T���|���y�I�p^�p��� 	G���n�I��m$/���({W�$���W�0ɘ���d������f�ad���Dr�7�5�?ڦ-��n>Vf@�܎�q߮�*tL��:b��{����X8���ӣ�	��V���>���1���kw��yc 3u��Ru�%n���PQfjC;'6����R:=1$y�Xu+p��k��2�W�l�U�1����<uahf�_ҳ�"�y$c�s��*��f��{�.#����zԮYj�]�;���p.a�h������|B?y�n���`0�z�~���F?N/�(�x4�e\�3*X�9b$@ �-�����N\}�QD�&��2�[ެX������X&�8����p[��h>6�˾��H�]�"h�Obθ�νFK2{��ꀝ�"ә������'K6��5O���k���S,`(�L�F�r�^$��!�>vAnEؖ���׬3��&9R�g;j�ɠ8�+?}z;�����^�Bg
���ZԅY��4����I��|�n9��/�х��ĨE��-��j��-��VSM ��SH�B�����!ђ��/��^5;`�Q���R���WF���q�R�E��u_����0�F2`bOc�00��]���p7�
��B҃0J�'�J�21�>L�oURl�X4�N
�]�ه����Q{�$'9x)��N1<�t�8����0�F����n]r YTy��<����k�a�*^��Z��������l��C_ü�H��4�^�`��) G/(2ljlVT����|�\g�_�=�c!PBxڏK�(�l�� t@�G���<��#yq��a���*����ieGF����D�d�h���`��҆(X.��D�esi�cw��ޡ�y�p���r35ۺ�ܟZD¤/`�]��yZrH�Y�ڶҴ��1#<�xoBQ�ӲK�\@����7n>�gS��v��������Z���C��j��WDA�`���_b��dT6uԫ1��	ܤ��m!]D�쁊a��4tL��F�.��~V�moZ@	���"��I�nrknVtSN��tԗg�Q�B��82%��˜��ҵ}Ԁ�]�=?f�}ޮ�}{�UT��y6W�U��J���!N{�u,*��ǁf�~��_:�an�
�)]�'}oy��7m�8��,�,���0ޫ� g:w�T�I�8�\����n�Fc�pi���'1)N�D�РMD�M:a���ze�����5�ǟ�gM�*�E��?�`��-���5
#	8�`ϐaP�}�D�y;_8u���!�eO�]��%�A�^v��y"�G�:��9#A�Kd����2�J��j0�ԣ�Y���x垱���7�׾o��i#O3�����M�-B2�)��'M$����r+[%��R���8M�������J+tZ�������?�H�ם��=��[73���"��htXL�o���U ���R^_�9= mS6<n8��7��;>Q����G�y��)�(Ƀ��O�^Q돩����c���HP�Al{�6o��# �"-fw�"�%Ԉ������S��!��7Q��Jp���k�p�h
�rx���'mKu�U���ѫUie��{��6��|�àc�?^�ɭ�D�5�E@��ǫc>��'�*���Qʬw@j�\��?+:G�\�W���}ⱌ�~E��|kI��9��j�=�Ď���߁W���s���*��9�Wn쟱�����B֨>H�p�=�����5У������x�	!��
���A>�a
�Asە�	x��"�q<5�Uw`	&9�ky�M��wO��:H��`���� >�*GwKH�=e��-��0y��*xq��8�}᤺��j�P-�������): D�X��+�{wYYBj���iV��q=s���Xd��~���3�Вs���
N������D�|�hK�S���1c�H�k��y�M_�N	/Bqw����M�A�cG2�G�xICiдA�R�U�*--����3�C�$kx�M41T8�)<֒�e޻�l����N�E�?��\�lR�x/��� 01�%ɮ��l�7%�� ���8�yC:=��^�)��o�D�V\�
�8u�{,?RB@�_AD�����&�W
H R\��7�I���k喑{��,s0h6����囁����Sc���J��c^��n�E�[��kh��]�ʐ�ؠ��1Hz��"!D������D�17(`U��Ly�+�E>l� �Y�S��%�}�&^�#W<��}�o��\MSDG+e��h��)W��.ˡyo�ZH��ym��?ST����/|��o�Ymk*`��	�B�9:)�������cf:��GM}	��8�N��O��6MF�puԌ'��Ļ>���s�<����,�k�UaO�qp�CH�3�W������*Ҫ���mV�Z���=��m�[�����	�S�C��Iĵ4A�����O����I��{�gQ�S�۱�ŖI	lԮU@��˭tc���K��%��ۥ��[����;�����Ĺ�\��f��M8���g�|�^׆�a�z-PR���_�W�����(�
�V�+�Z^L���8!�����Ą�M�1qqL	�[F���M�HY���7��Ӟ�ˮ,��w+T39l��-����Q8�(4p��e��PF�-l�{� �
�p���2�&��L!�m���c-=�i�U�(�v�@0Bm�>Z���q@�g YDQ9ȫ���[�.�v)7��U��3
˭�.�L;�����xJ2l�l@d#�C,�"pD9C2 �c�E�
���&�&��n6�V�Lg#��F�~[�zV���詭�y��r��|	��K�M�8L��뷚�$D��9gѿ�,1��#���\�)	����`2�rn��e���y3ܶU�@��4���F�`�>���غ��W�B���@���r�#�z�����/�f��ly|dbB6��//n(k�+N�b$�i+㠁^g=�.�vH}�D_��jxZ헥(����"H߂�d^�I����P�BK�!�g��7eVB�B��M�}�����ux�����w�,����1���L��%���5����&И�5��4�Q^����T�(BF2��ղ�k����ɾ/�01'*�q�Q~�>�����l���/Nnd�B|�%��%?DI-*Q���&D�7J۹ZD�?^���@�UdN���/����23�R�y���x�6��z}s��7}%��J�'T�|�i�]�*AD�	�=<>�r�*=��v ��<�!%�j�F�xe�\欗��_ � 4$�/p<FZ��5VF
3 �J���:�ޢ� I��/ �Z�K�QR�a�m����C�z��!Y�3����ĥo�U/�[\�1`K�"}�Ls�!4z@C��'�WG����7 �l�q�E=f oN��b���|����Hi	�?�P�}N�a��p~xO�Klqz���#�0���{(^x���Z4t�ؖ��Og�Y��jwQN��%��7S���vaz*�A3�Rb�Q�Y�
v��]��8���.��V��o�B$��:]�h6������zyr�CI,M+����nD��I�|_�r�WQ{*�Ĵh}�O)�L���eՌ0ꬃ3�O
���"�i��'ʔ���K�"�,l����={��7 �k��~�w�+����ޏ˓����g���e=��i��n�+g�T'٧��kV6���U���>�|Asu�?s��/C#�Hf�qU����~��;�E�&rN�/���
����r�?����tc���gqf��<�/*ޘ��Id^LSC���,|��@�XÓ�w�#��>�f������F��t��+Z|��VI�=%���6�ˣ�`3��+pD�m�C�;NWuJ�ĥx�F�V✔��6�	Y���c�;>ʽ�`��ت�&�s�����5��o����{���u�ѕw�p~t�_,�AW�}��}��L���e��$LoV���X�o���$⼀��YX>ɒ�ͤB��")f5껒R�q�����	k[��dF��|�<uS-R� )C2s��Ȃ�}R>ntPŁۍ�=*"^�UݮwԮ�������n�9'i�L�@�Ǹ�\ON�deuz���O	I.���7 �}T�]�bǒ�E�Zs����-���^�y��N:O����5	����g�r%0�q�aW����CL4����7a�ܴ�5�헲X��2'rlX
��S�]��R������[]Z��o����Kw@��'�<v׷�ڴ39�.hS�����ι��=d����6���G)���| �*@��*h�^�L\���:9~W|��b;'ǂH8�K�A<\��Ws&o�J_1�`�����Ii�<�"�:z�eXwo>��u�RZ��#���W3 rJF5���^ŕմ���'��-S��q�{�؂��j?o�V��Cq�߫��ns���r�5s7?��(@�t����m�Jo_不l�n|%р�.�F���LG-���{�N�%̘��:@��3��ô!*���i�O^��G7�ߕx�c�f�S���8�	��3)��J��lU���PN)�x�� ����4!��n��������
I�]��U���s>�*������8� ��"��aQ�����tJ�X�����#E�"���
'���
뙺3�#9��\J=�K�s�Gtw+"l�y�Z��
��nYN�	�Z�����`���̚��@����W�kkUcQ��Bߧ��\�v�~�
�������P�Ь~/�f��f����u���1���S�DY�W����j;�XTS�o�fA-����S�HY�W�*�ٳ!+�ϑ����K?��]7Wn��}�q��qu�i�ؼ�� "�]�d�� ���8��iޛ8'�������ٛ�֮D���v��BA�҆��6��ooM�ʹ�-�D�f��E�5���<TZ�^�x�@�ŭ��7�
�]<�f�;���[U�i���'ڨ�˰�f*"R'��L1!�t��y^��@D��J�=F�_s����!ܕ��$˶*�p�gz�Mc�qE�3�o%K�x��`����̒�U$nFsǵz̶�{�+-	��6}�L���)���l��� e@�9���A�����5z_��^i��4@T�À�t�C07�qBIc����`4{E+�\�j��ߖ��(�3�KtM��P�$$��.����&�x�o�i���M���"m��������i ,��c��@�H6V��SϢ�:�d�F�f�3�2�h(� �@^"��K���ԓ���c�6��4D�YM�hz���-���a����94��}�)�~ȃ���ƈF�+��l��c�RB���V���k��ĥ�a�����ɓ�W� -G��	 �X�MFz����ZU-�$��]1���hf�\����沿(wYpM�l��θS���C|�|��x���z �]�͍���}"�2[}'ɮ�6��+�N\%�tzŇ:$1�m`�Ê�}�ZNj�H��\�еf���"�bU U����v7��t�y�v|X8�����n�ɗ*V���l��],h�@��K��Ca���R�;>M�����n�E���o=h8�����@�T}M����:hX��!t~$�o��YiÉOP�bŌa��bA�4�k+�m20�Ι!Æ����]�a�T��Y�R� �zz����eɘ�����4ϡ��r���j+ol��[�BX�����2+��L��m�n�K�w��)=�ϗ"e���W^&��4��	r�ƣ(��H��P|e�)T��%r	��(H��9e�F\�tu���y<tw��s�����	�ɅN��qC� ��˙;|~�<N� �?�̓�����6SߎZ���?����>�LT%q)�ќe�؟>���Pw�N�K�����>�T06�|-�v���K��Y���s�<*�dcO��zR�-͍믆�ع����o�G����&��ц�y���`�>X%�ixd'�M��Xdk��6h�(��w֗��u��L��������{�mZ4
�×����?_߈8�M(I���dɉ�Xn��C�C�.�3�e(��C%@#e�,k��O��!���&�]+�i���H�&C�剥w�b��]D�R/N����r��`-���{�#}���.�²N�?.D.�V �+XRz���S�6�c9io�tuKP��]ե�V5M P�r����&\KIz�)���Z�N��s~�<�I�\���+�;3�����n��szs6G�t;-��g.)t2���|kP�e�\t�7�6w<��M��鋡���&�=��jKV�c�F��
'O�ǻܨZy^0�vC �����[ٗ�+�öϮ�K]su��$b0�|��T��n0�#�
�h��IѲ2[�������@�aiy�z�n
����M}�sb\�=
��|��x=
�I��1kPIhg޻���IK��D�J)7	��y��'�ig��|+�d��y���S*}E���ص�JB���u�|d[�L9L>��3S�!m��v�3?�N��O	�z;$	�t��.��-V��`ٯ���eHk�I�1Y�:��S�f��_�U��í�)�!�>{!�$K#C�p"^FڎBt ����x����^ӈD�̿𔷴p/�
�SpL�N7`���Ƣ�@ޕ&�KP(J5$��A���t��i (�Kي�S����c���ե�Fwr��քJ�Hw��� ��B+��u';�"�B���U�� ��'Z	i���+��JS}�%~�03oȞ�����g��k 9�Eݥ�������M��)NI��"�W�^��ީѣ��vb0��ؿ*��ga����Vɷ㲼]�g��H��M8Dl{�<P ��iZ� �Pa�l��P���ja��_���Ȯ�������������ӌ	�/��+S��H�`����-fL�{���ג���Zv�*T����h�ƃ��&�.���h��g�R���z�	.k��au�\�j���g+�{� �a�L���L�#wB�L��:�y:�4�Q�\D``~T�*�}��9+�a�NKH�ߒ܄ģ��}�B:�6>����^/�9��ň}�zQ�����sr1I!��+h��!�E���}h	pj�ُ��V2�`Љ�<�}r�B�a�/��@�+����n[P�句Rh������}�r�@��u���W���{���1.0�d��PxJ�kV\�a��w��Ax$F�_�� k���o�9QҌ��RYdA��J�#6�tDX)�"6 <  ��+�+�T��X�v�W�^�������m�{���l+��jI��jc��jf����FV��Џ�q}!���� w��c
�f���h©�uL�eq��h�aGjT]>7��`)�U���
t��h��7��F.a��L�a n��22Oc|�r箛�c��Q��3�+M��
l��n�:o.�@����Z�u�g!��ɮ;G����sU�B�Dw;��\�vP5�]�+�ᬶ�6�6�3 xЎ�O?��Dvi��A`h��!�(5<5~��Q/,�
g��Oȕ�e,�?�L�>+BW
gw�S����ep�P�^+�M��� �p��F��˟�c�M��G���������t�z�o $��Ǩ��.ja���6���f��ؾ�ȜM3h��[ȭ���B�֯>l�T��o�b�d =�Og-�L�֍Z�ؙ�#'+˂�L�pܥ͒!�"�OR��;��O�\��(P�T�&�<� 7.��v���ʏ��f�B�f�HO���X/��
�% 5ń(l��fj�aVb�"�s��HƤ��]���is��3p���->��s3���P10�r?�'�Ė�p�J��������� �
:JI���N_DU���ώ٦��S7h�_T�'��	�l985��م��*{��"p��6TP�9Õ�Ŗl����G�4���|_�0�C����e]�9�I*tk��S����d�UD�G
��U���n�K2/�D�oB�vb��qKz���E��4�Rȴ�f"=u4�M�X�����:\e�G�5zG�$�U�#�E�x� 8�s�������<#�,�Hn^��g��7��/�!�leҝ�	fm\�s��+��:k|-���< �퍆�ؗ���6���C}���r�G��ɟZ��P�����l��u
�X��챷����N:�j��=�:��;�5E��r@��]&��>��Ә�c��k����̭R�L�ג�&�Tꢫ@2�̡�-��wL��DEnɵVU���N �7�Y���b]���v)��H�|$8�;�<�\{+��%�%���"%�Dڬ5CwY}YېO�YT�>z�&i�an��O�G�ـ\���/BȰ/�[&4ꞯ˂p��@X�p���ʊ>�.z'/�0|k}^��Sp�(��S�ʤ=W��L�O��µ�A��k���,J*i�"��##�v�%�6�B�q�b78�4���O������F�־�/��c���'C rdTh�&��FDkDW��Ly)�ݏ��0�5��j�F`����{����A�*0ـZLȖ&W���p*�_tK�r�R፬ǘ�m���*h�#Zi�	�(�3��5�����={��m����$������\`YO��$඄+B'D]�1�E�����
�5`:!ex�2��btT/���NYexB��Y)�*��#]
S��˰���Ȋ��X����8e��(ѢS1r�m0�cp���h2��C�O���4$���L���aۛ�т{��+���r��Ő5�`ٿskC�O
0-���mo(��+�MK-��7Q�!��5��Q-��5�2]Tg�4Y��;2�����<������D�26ҟ��U������J� �:��oRw�zC�79 �*Z�-�(Q�>�F��q�P�&����Q��svp��ڑ$��6$��>�C�x/�s`9X{�Z��!Q����,�������]��0�r���Q�����J���}�M�nmҥP :��S����ł"�~���֋ ZJM7�T�7��A-x�:�=v%�-�M�)[�l`�bt�IWI}��x)������o0�s-�d2�Pf���hW/��2'i����J�,�K�Xح<)^{���(�z猸Tt&��FO�d��h�
���j������_ꋛ������l���Лs���b@�ĩS��*-x�t��!�9`�+��\��]HU������K�/w8��W,�S�pT�iHl�nÉ
��������s��H���F\ő�����4��D�g	�n[��8Q��I@V\��I!��V�"�6��`�lB9$���自yqP���&��픞��-*\�\,� �]:|\3����Q˒XE��SO9�1�iխf����:ՈZ����aݸ���ӦC�?.ed�>[��R�����,#	AG3o� �!��&�I���m�O?�ۜ%��˜!��"�8g5�j�ub`4�J9)���'��U�'��2��E�(V�ʐ�t���9��|�]��^��
G5�Rpo�\rP��uwē]�Qgͣ�W;�]��"��{�
����)�N�����L���f�����S��&��1�rM�ݠ�KI����6�������䔓�:2�����������?9fƣ�hE<�T��kR��b�-�3��H�*ɪm�B�,][ʒ/V���c���>Y-�L�L�����Z��v�ȥ��l��I��=n���k��@�e�~�ĵ`:���-m+���B���۶F�{e��{�˻Qݔ�0�1�����ž�>��K*6��)(����W���y���#�>ef��B�nڐ�=�1�9�+d��-Q5�I�P6,�|b���}�pO��-m����k�ً�c\�6�G�9�4s�P6�S�K̓:���o�9��w�Н��d��5������eg`{��X�R���ӧ�����"+�$��)b)�܃�*���f�g�t�#4�ʹgim�B�=�+E��lP����AC��ˊ+���8�];f���wǢ�� �)�IK������^B��	���"n�\���B3u��c����T�@/Hk��)t���]6�da�^0�O`o�M��V'"AR�n��գ}M�Fp���u���|]�~�����'�s|�y<1�Du��ǘ5�2���
O[���aٌJX�yXZ;%��#�8�-޵��Jia�lq� ��_�����^Z�������I���n.ńD�����
��c�h�*ZN�{I�S�R�o6�b3�>�Yм�7�o��ܼ�ǜ[��|$L�_���_%�/��6ul��E�1��%t�dW6�jAPl�g��(�A�zxy�Nbޑ�V�*�s��$�oc�=�O��{3�po��z� ��=Cq�1�z�C����m�aǞ����
� f$q��YËXI���wU���_8� 4w��B����	�WI,�C����.����HR�tDj�;+���x~�1�j2Qi:�Kϑ=A�g�ޤ���F���HetG�9����s�i�+v�i�2T�w�n�����ݻjx��L_�\�b��a ��\*X�(Yd��I:�V1Fq�1s1gK�e��fk���w��:.�"����-�������ҘsRS�¤�7u|�8��z 3|���)�[h�kW�%ϑ�����Z����[��,�����%,s�T���P��}��XH	�2�,!Y�@#�$�7�q����ÿ�<���(4��h�����?o?DbCg�~bL��q��{%�,�z�?ro�,VIX��<y��ˣ}N�5�p�U9��P��dT_�3s?�*s�,P�v�?��Ph�#@����g���=�w���9ƃ�����:1��Gg�f�.en��uh��Qܕ�������(�iRi��N��Wӱ��E�{|���롬`\U���E}!/YK��Vl�rv��pR��,�6�1��q�*�S@xB���,2�]�4��}03P�̿}��ƶ���o���v���(��$5ɹ�L�/�(�zg���#�:TH$d�)�#
�������+J>�DD�u����ߣ���d��k2x _�)ɘ��D[�ku^���2�E ��C�Al� �ܮj��&��xB�j�SR��)r4����꿊���rb&w�4[�m�F=�k`���F 䟓�=�\�f?&��o��]@�p���*�3�Nr��O����UT<���9f~����ćU��O�{d�C����D����^k�}2[a�D�B�iI�OS�B,���6�����4Ă_�i�!N���?B���1t�˷�"��X�#(Ӧ5/L�L���x]
s�N|����)���#m�`}�=�&C��:����_,ϼ8��r*->!�A��K֖A�i�(- ��[�2d�\����Q�ގA�<���a�$��z�����d�����,�|��^�[����}����ט�S1
��z����>��Kɍ��JD�5���)q�qv����Uv�8fN7�pp���#�\!9��C�
U�y��<� �}�f���7M�T��Bߤ���+t�V��~�*i���D^Ig��$ʇZ;>��}س������l�S� �	��~�E�:���#���(�C�3巏g�v`�g�T\��60!��"�}U|#��,�i����p~��Z��F�U�`��� si�l��g��oܩk5���^5<���$ȕ\�;�k�x�(�~x)R*y�.=G4V�G��T����[ς�R�k�z%�^<��̾忔U����[�094��/�Ԥ���ʕ�R��ciwZ�Q��`����b��@
{�qm@R�\k	W�(��3�Z](���3�t�v�J��?���>kƙ����#����%�������ZJ�6b�jD]�b�U��P̱����&T��#�o��=�eC��?ϯ|>7�g���Y)}��*Ă��qX@1���'<2�5g,�.���4��ՙ���lC깩w�^�6L��	�y�~��CYaI�$�t�9(E���y�y-F�� `��Q�_������e�r�q �����K�a$��of�eQ��Oc����<�J��%E�a[��}π`!�}��.ˎk��ltF�,��`���i��/��4�z�DzZ�����ؒP����-R�q��ճ�W*%�$T�g�1��"����G��I���;(�����Ŝ�8!��BW�&갱�
_�r��%��P��ٲpw�6�$��o%�4��ޞ�f��BA���X��Ls}��"�y���iS��c���'�|���o�8��X�1/��N5���QN�a�������|�j���(�L���Q�B{b�Gέ�${���w<>G֏��Ybq�qv����=-��|�f�_'��D������{iB4ճ_W���f�L��Q8�<�*hI���m�kH�.8��c��kŏ`-�	��ݢ�!�h~&�iK�;S�*!�xKYz��i�NQ8ɹ2%�!�"�BkEe�D��ܶ�i�b72�������*��ŋs�ƺ�.���EZqs#�Nb ʅZ��'���}?&�ܫ� l����?�2� �6�����}Y	^j,�����}�ܐ[�^z�p�P*�@�)��N֏�(�?�b�~ֵ�Iq7��!5ס)��y��9g
�H��[�dlIL�$~�V �|�d���8LI����ަ�'��m6�U'�uk��Dط�ʠ��q��{R���5_
�U��e��[A�iO)dY��f�S�b�+�q����$��JC�; ~֤�GxQ�I�i����|����-5�"�tN�C�u(�w��%���f8$�}�
�"xj��Qb$���h��ЄL
��I��0�� ȉՁ'��^ͦ�D%�J�?�A�D�t?u�I2A��dB^ ���c���O@(T����<4��;c�m�R�����UG���eJ�]
���S����C-ؾH
��ȳ��a'��Ů;���&������w��I!0d�_)��pp,GV�f�X(D��	����Q�ש��|��g3IaJ�՘�i�8w.�Zn�L�� ^K�j���r�fL���wA��L,��BP�4[�uv{���!��FZ�ډ�JS��̮
�dB>H�Hۇ^�����"G�$��c�M_V�^�z�}��ATs��[�*����:m�	��p�/�>\�17����R���w�He�vn��O+�e

�\�GhP
�����wKJ8�f�:iP��vjfyIx����G/��׸��I�a��'��F������'��@ Ml����`�����cjp�G�|���.˅c�-��L<�gӊ�}�ŞOR�Fm�c'�]|y�yåE)7��j.Ť��w:O�hk��DJ5:��USn��"����\�H���@kF����.�5�1.`���oa�$�?�	��ĥ��I~h��K�4�ȁ�a�]��^n�7�����������к�Wt��N� ~�s�	T}�
�H��G|��$ '��_R�ۦKk�VgA��ȅ!X짥�����{FAM�k��Ţ8���M{��W0pSC��4cGO��d�M9��m��zj?�-"�S�+|��Qs�߭���Y��Y���A�N;kL1���`߈�pIvف��Cƈ?�����t�I���&	fl�=�uX ��3s����bg��~|YFꡇb+!�|�������������:M���߸�YgWI
�1�򚟮��s� *��D����`W��VC��A(��*t�t^��Q�OM*2W� �XY���F���?��I�2v=|V���.���.P3���3�bL�iE����#e4�F�N[ӱ��]���<���o#�R���?BG�<M��h�1ʍ_�'��k�0�L c�.��vj�tא]~�	��y��=h��`����ά�n�:V[�������P̠�%�`[e�E�g�H^�.�4f(�?����Vvd��M�+K-�@Luʼ����..�_t���2i�|��3'�E�F#sitXs ��:J�,�\0Ǣe�(O�>���>z�J��wJ����[��!.L�;-�s�$D��|�_�xX�f+���+����o�#�$A�:+�]��X8��IP0{76,]����_c����yQ
�US�$Z�Z�yƹ��1Y�������J�5ޝ�3��W%�>�Qޕ�7'��1��behʳUo��B���l	���Ҷ[�U/��;v`�'e��:+�m�Q�J��7tY�w{��/p`����	W	�)ʋ�O�1Kظf�|��f{��v�j%-��lsX	yn�,�Ϲ)�<���e%6�m������Mv�Vtn^$�H�	���|��KԵ��[��ـ�E,
sp�݌���-���gf�(:4	}d���b�iwno �~��u 7!��*�7�v���Jq��Ȩ�5cr:�6Sn8�lИ�XC�����'S��q�b۫��P�CsQE)g?��	{�|vzQln��p
�^<B��b`���3�!0�~>�p���s%ڸf��;�S��,y㧮d�H��Ei��Y�"���+g����#uY1<���/�'O],܄L�3I'�Y#�9B�8�c���5�M&ʭ	��ɭ�b��S���)��C����it~U�����~9�a�j�U;k��d�s�{�h��l㓢d��*؜�$D�8�����9�J���-R���mع�L�+a9�ap.�4Ȏ��z�0�v;��7�n3�XL�q/�|��	��Ө6���X/���)��V�M0�Wɽ�j�%���+����On^���֋ǂd���4˥q��zPV�tE�4.uh=DaI(g�]i���o;m��959���1��o�e K��8������3%���1��<Sc�7��m�d��#��/7���c�=�3xQ��ݏq��w�̩e����25�դ�_'�'\���'+�<m%2�����c�r�z�*ҕG��a�So���r0�@)rޣ��gz��gXK��P�Ңd�=����,#(�T��F�$�'���\	!�-����e�@�jaUE�U��P!��/S����o�p�底g:d��A�4hi��F�z���@�i��荲>Ēx9e�4.���u�f�.]��qk}�pN�*H�i�ˈ1N�Z6Ͱ|��cj����{jJ���?�g?��qN����Ag+�K�T��*Q0Bp�NA ����!L���������A��[��9xLVD���6�����S��]R|:t3�a�BYds*�oyzB1�GZ��!�ukk���4m��_؅v�ֲ�-��c�]�3ep�HgV�$���*Y���8��Ly�}��Y�@[��܈@��E�2	�ۈ�-�2W����bڏ�B?���c����0G٠s��	�9�̚t���W��y2��zېd��ny�U�����v8�`	��1?�͟���3��2^�h[�D���B�
��c���ޅ�]���h�d�&�ǔ���8f��~� 4�Ǆ��?��K���>��Z]��u��a��u��_��ɞ�!QS�zDg0��#��q�@�Ƨ�ժD%@��i��p�S:Z��-a�	������V1�Em�/q�D�x=������`i*������H���Tՙ������<��M)�-�ʢ������������Ln�렱1˼
u����!A�[��Y�\����!�<3y�*Dw 5�C@�T�V��3ئ�T�s�e�_�\m�YƯ=���l� (�`��3�ڒK�MЙ;�lZ_��9���6�Bt��Tqp��{�>w�^oN�c�̲��ѷH�r}%j�P�Y�י��fσo8n��{�FR��q�>h�t䴃�(���~(����\Z����\�+�K���\��7����?vs���Z�:���l��b�������jmG}���j��Lb1�"�Q2+Gʸ���-�b�{m=�	cd���.?�O)�Jx^0%ŧh�-ZRu�oW8�s��$�J]4>��?��nWc�ϕ���!�F����!��� �S]�O�0������׆�ZE��U�������g�a��}���$�c�u��5���H^\�������4Xڣ�Q�X�����^{�~�^S2��q�'��X!���
��� Y�{��H$<��D����f?�_�E��0���n]@��21��,]�P��?b��_��.U�����1dn)�hs����E�u0�
�`��oI�0��)�mtzJ�{E��J�p��6�p")��F�&�G|ju�����O�R3��W���#����m/�r� !�cQY��ٶ�C$�8����JT&����Z~;*�i3�fH�Y��)�4�mF<;6�%� �4OU��w�9ߟ��郹 �|���/��� �-4� h+��su#��Ǵ�5:��AL�J�yaI�P��j���_ZU�o!�R��l7YܑX�)�".
����ty`
��:�hfG�!v-�o)�Ź��N�hq8d��P����ݓ����`����Z��&�)�Z�ʘE�9�k�H 1I�Q7.^X�������f$��h�U+;K��&\�a� �	�!�s&�h/�qcy�-=�Q�Af������V��=IW�wnM�����qW�t����]
��(N��U�1�pL7��ʲ-l�M������ k�~�X��K&k��I��]aKM7�t�+�4�z�,�OrG�3��_@t0��rM����xA�@sȅ�ۈjm1,�,m�-z�����}<Z��Z|р�_�e-#��N
��,����3��3I��蛡�$٢�$jƳnS���bT.ը��=f�[T��-<չXѡ,�5��E��;Ɵ���W��3�|*D֞�=�̛����.ŏ�9��k�Y����T]Fe�X~wJ~����&Y���ބ���.F�d�H]d��!�V�U�$_r`�>`��e�w�ȑ��K�����=>���.!�ւ�V��t��\k^��鲅�(�48���9�sbХ��tH��b7�z}bzx���#�_(T+�nX�e����WL�G:��4��|'���\�-؊��Gm��3}q9�XҪ�:0��"�~Η�N���+Xx���AbL;+Ӗ�rA�ʋDϱO���L%�ݖ9�~�h����&QU<I*�3� ŉXf���m�A�N�w��6B_��?�)T����4��a��"1c������z�-]m�sl5�D�u�\�_wU�������x BkV54F9�Ab��F9�d�1?��2���*��C|��oў*����������C>����ٵ�l��G��7I�w��f{��~��~ԅX�������73��E��|�����[[% i�<���U��f�W����n徉�%%%�H#x0���]��\�᳽��4n���i4���}�r��lV,��L�ot�?\����Pˮ)�ؚ�� :�L����Cx���k�%>�K�۱2�z,Ʃr���:�G� ��:�Ñ)pz�Px��{f}W
d���l�=h��6�\p�o[ᚡ��\��E.q1���~�W��	���y����x>�_I��k�6�82��/���8�v���]�<ko�H_2�����.4��e���&q}��},�kܵ��4�_v�2��[��z�ύ�gd�p�߶�Q�.���\�H�1�u3"�pm�(�/QkP�h��w[-n���W`�#�q�a3�%��G���sq�R�s9wr��!v�`�Bz˕%��+���Z)�3�	#V�7e��{������!U֑2
 ��B������"՗.b�&�����[=r��`
a��!zG#���s�<��獤��u%�4�8���j��k���l��.�|g������r��5mZ�e���t=e��"�o�$=�t��hN�"b[]"+�"���z����x=Y� h��W�-��D��g ���+�� ���1�R�ê��tv���L�r�FS����y
t(T��}q<��X�F��ЕR�d�N���~]�j��C�G�����#�<�x�ry`�ᣓN�s#:^㝌>����!�!A�����S�E���x��w���b.P���t��D=��48�#1 >�:�Urf�c���� ��rl���寳�5"S�"����!f���©ak{��(��>W�l#��w#q�����в�?�'s��:�?�Џ��2#ꂱ�5-)�Ox�3��p�n�����s��Yn�r)�����Ɯ�j$I�_U_�,�q��͒�C����$m�⭨D�\,nq_�DF��ą(b[��2������ds�}������S�Y��ϡ&��s�#���i�G�ö.��0���d�[�)<޶�^ *��pTZ���e��������G����R�$�{�2��N�&�|>WW��8�3��I?檙8Pb��o�J~L,�rhC�VSl$Uh|U�2��.dsZVa��eN�<M��q!O����aġ�#UNWb\S?�U�fID�p�
���>��K}۲6:T��ȱB{Y�ɺ��;d!���k����B���g(-;���c����L�`��=@��l[<]汪q$���.�Ac3� D`�I���*lU߯83�;h���˟�U��x�Y�b�)�׈�5�V`?8�Ԛ#��Ԥ�iˍ��6��'��/�w�K}� F�$��[P��f����s(ZpK�u[Zsg۰L풃/�!����Lb>��	�Vnŭ�"� }���O�6�L�#[]İ0{����_�S&�d�?��T_�\ί�9PpfO�g�L��A����c�#l�"媠ha6��~����������?f�1F}0 �O���4#���Wp1����<Q�iv� K�yAi��G�#U7�3��Jj�]2.g���p��%ߟG_��vS�VT漝%|��LWt�;�#�m���Ӑ�젻��A�ܿ���uI�>���m�]���V��p�sX�&� K� FHv�7d��\qj���;���`چ����EJI�Տ�U],TP��>e4�c����\2žu �0���w[����F'3�/�!{�������Oh�
�ǲ���b;";�UsԲF9����ھ���
�t�^䚭�[�+���2��٧��l�h��Z�>���C���f���N���*ND޺!�"`�������^}�n��;�*��ŷ���a�ӑ�iu_f�#�=0��2�x���W����H� D�Cd��4,I`���b�i|�����cL�.=�o- �HB&�.���A$�fY03h X�b:�ј��Va���رyOh�y3�sߎScUVZK�H
vl�I���+�+j��tO�H�OG�n��|��Gtvp̄��Q��.�ɤtu��X[��*�I��/��V23��L��u�ۃ�����UT��2B�[�	zr�Br��h��i9���փ�����53$E�>N��BIl|ԩ�����a���2��~s�tG����L��%�|����Y�Z�6_�c�M��5��f�
�C�����!g��5���Kv�]U��s��/*�Y�.<�bG��n�P7 ����R*�0�e��R$�\���:�|��d��X`�&�a`ڱ�?3g��K7��K`h��ݚ5�[��X|�LZ�6K�33��Ԧ�+���s2��i�/��qp\z�A%=��y!d�M��2|�Z�<���pp�uRk�~�_,�OZ|xJ�'��_�#�%b8h>�X� ��������%Yu�^>J_(�u�Wk�ihI������$u�;h�1K�d�l\���+F�J04�9}T�ٴ�\�2?��5�"J�u��ۍ�Dx����~k�äE���aʢ�-=>S��P2�&e�!��0����7��TǬY�\.D��b߳��D��8���g���>_�y$�y4cD�#a,+��H�ʿ��[�G��6�TW��H�Tgc�7#����6��f�M��,[0�rc|�U&X0�	Vqp�K�w ]$6��;�z /��[�6�M� A�XV LO7>�|�ܰ�P��ᬶ[�/7ܠ���w��;�r�Q3�NX��K���v=�*���-�`�o&��QT�)Z^aҝ%���1��9o���V�e�0�E!�Ϲ\����a��? {�@!�����I��0�:��C��+L�!�fI�Z�������> #�B�%wʉK����Sw)��RK{k9��)�8�Z2���i�`�J�l�Ԧ}�=���n1�K/Yi�E��� k g�z%l�}� �Cl����(7����H��U��ݷ��"�.?�s`9�kb�����m%)���A�Na�^��#��ٶp,��'U�C�������QhS�������h�\@���gꊣ��8�(J~͏"B�E��}TYy(�IUD�(w����)a��L{w�r[��3^��%(Yɕ���y����Swcr�Y�����_�F�E� J@b-rO�j�\b7XI��jZ� _�{�^�
�3Yv��_@��5�ڮ`ڭ�[��#ńa���t_#Dȹ�c�A�t�d>�A��r� <(����U�x���X#�/�\uYcs礟��g��VRXֺ��������,=
'�!<&weC�`	ͲR���ϗ�u%��m?\_uTzϤTE<�v���zh���?�:�_"쿫��C��ͱnq��0f�i�`�bE�3m����;�W�9����'E�tgB���ؒ.�E��T�{nz���a���h$���:��~���P�����3X��µJ?܃]��G:Dİ�.V�{)^��r�{�l��q������w����GQ�*��F�WKط��"��oн��rmӷ�s/*��nqnc�cА����Y�%>&)�s(F|A�^,.x��)��1J䜬�m��$*�v,`�q�?��zS"bt��M�ĸA8���@�P �Y̷��������'�qG.�"�T�����>�	���#
9��!�K�H�5.%/ی�L�� û�X��a���8G#3vzb�\���kAl��I�SS�O�b�4{�=�c�Z�a��(����l�+��i�%l��*�ƕ3,(+��T.X�}�yޒ��p.�w�QE�����iL�x'F�-V��δhZv�����0G315�/�����FB����n���(T�Gf�0B
9�o���K�Z�n5��8*�������]��9���m(W�P9*<��-r�X�R;�dRP���!T�����x�����)�d��/���z^[�^j�b���,MI��4	2���)�4�!�Ӫ��up�;-mԥ-�D�p<vy���;.�u�Z ���h���k�#4@-�D�U�C����5��W^
�Sq�∗�t?��s<����� ��[V�@(8R��x�'NH8/�^�E�|Y�0v9�1�I��d3�Ę�:�avOjq�� =Q�rm���/D���ſ3�!��=}|�����ЯF��X��9l�7��r�T���Ӷ�az�����DjM����}����yP�5y�#,ת05��U"�a=[o���6���Cf�#��Ue!#��&_	�ȭ�t���Z��y́;,~lt���O�W�.4���oI�w��=��������s�
 ��m�.
5��Tc��B��x��J��"��T�^u$*eW���.�%��.xg�H[��9�G�#�P;�|(�ؐ7
#��Ӭ��3���n(~�M�adz�_�G��lL�y5�$3\l���'j��yJJR:�
�34�.5d�J�4�̠r�0#5�U{ö�t�0"���Q��˺�/D��e:
�A�C ��l]$��	ʪ*�@q�Pխ�Q}X����n�K��H�.����7���m����������.$>��2&S:�����p)��q�7��u3SH�>5�xc%��a�|�� z�L0F��������l��v�1�Y��qU&��������Qfg��� ��<pX�]����d1�G�>��M*����J���Y:�iK~r.�G����lQ���H�*��l�<���x��9�my�ՎLX,�a�#��`w^�����9q��?���|B�4��v����ʈ%�d�BX?L5 �N���L|H�{� 3%Q�І璉�<�y��,4�;`�!�w\��q��+���2#��o<�g����	�gK�c�ľ���	���\�Q�(b�$�w�K�Vx���ڏ�J־z��?�
)�[��҃1�A���� ���kh�̸9�UT�=�`�� (�-D"q�-
���M`1�� ��KI#��K����p#���Di.��x��.��[2�7��Vt7I����ma����w#��`�v˽�i�M�A�~�;��îv��7+ȯ�Յ�;��"	_��%�=>������/F�C(����5qn�LX�p��h#�3㛴�o�r�ЭE4K��� `p.�çD_�%&�na�dˎ����@Q�W�/���pO)�=���(K����y":@��Ջh���*T���{zه0�Q���	R��\�5ػ���ԛ�C0|���>{N{Ĝ���풋�@]��|d�Bx+n��z�~�]�*D�(RL�f���.ݠ���r-��
-P����H�r�,��´��ı��s�yw.��jK]	o�OG%`��T�����Th�P��`�#�e���i,6�`�_�`+E�J ��|�-8zݟ%Z	%A��)�����+e�;.ҟc����$�*��E0hc��z�U�����'g5�p�
�\�B�1��:e�x�9b�P2h\�;	}{:��of�����3zT���h'Y���n=eJc�8�6bS����J�vX;ed:�	�˯�z@� p�͟�K�g��@�M���L���6�T��nY�=Rd#`~� ��Ϝ�S>���	k���x``�e
^=���}ٸf��#>��I�L�Ｄ$� ��o�ajejR��t ���I�n�+����?�7�̇L���e�dG�>� ZE)��6�����CݟI1�ı���ƿz� J�e��_S�`^	B(��D'ǝ�2�]P��J<D}a) p���$'����z�OT"δEJT�y%�*��n�����;�n�&u����є�VF�E�E��&8�¸���J�P^�|\�v�Q�K<�rd:~b/'���۱�18�z]��\?��~�Y��77�߰�2�<� y��a&��8����ة� ��%:��H��������s)$���x�s�u@]H_t͊�`����h��g��%�	zT�ws��(�G�0A�p��Η,ɘ�����4���I�Z����(�].��tF;LW�ku׉k�O��8��?=~\�$#�n_^A�vb��J��I��%86c��m����0�zꊧo�_?0�V�z̬��,������U�|@�,V5G1�y(TGz����b%!��W�ݒ���N�)\�6
�"�6��1�(�T���6e���݌�����u������mE��'����`��}?�{���'�A��+'V�۠H4��s��<�9@��ͺ(�1�[1�z[��~�J%]����B�
L0���1ڷ�a���ê�� 8��)bl�_�A�{fN��Jq��}_ݭ�?V���6�a�^��)(�'V�`���d���[f���Y�Z�"NEΌ�L��p7��s�u�n��8��/�*���A�uث�	�u���������A��Qoi���<������t��k�MC�0��?�1cǆH�٤k�N�1�W.J�<��_��	M����C6#A�/�7��8���3/:�������a���Aw��-k�	�9Ƃ��C�!�G;�}0�(�#�}��׆%��_�:T����Pl%5��E�F���)�d/n�ؾ�~8��=6��+�g�~�Ms��-R64�������5[j��s2~����߮��"�&�=�6!�O�U���渐^s����]g&.�́E�$�tp�}+�(=�Ns�zסTRo�!V�3���]�OQ�"
��Q?�f��[�q�q2����?)�m�eO�{�RM��	XpF�D�YB�s�B��҉C��/��?����N.$b0 l��y�R�F���$'Q|�A�n�E�;Ҥ��1��DQ[��<&��\+e�|i�v��%8L)5�8�}��an��������4�3���M��HC�c39�ʃ���1�ZY<3��/��N�j�}f�#Iٵ�%XM,�P�BP��
-��i�8�(�1β<8�7����mSG��
ZL��g�x��(_�R�$���YV�`׼s�CC��J�8W��h�uΒ.��w�T�����ҳ��?�u$CnaJ*	�#��iͦ�9���"��`�^7/P�3?>ʖM!�� ڧ���O�>x�="*LV�]<���]�h�Z�d咯��S�X�ww��p5��h�C� �zݯ{�Q��@Hc�X���r������	wv@1jŚ1L�kwa<��K�m4<��Vl��V� D��Ȧt�8��_:}_� \7^te@��6#��B�^���C��w.�l)��:��U�,i����u�/</�����7�o��+-��U�s���QO@��Oi_��ٰo�r��uD�K���:����� Y��nm�O�����11�9�m���>y
��1�-wpBc|b���7� �jwi$�6���
I�ξc���-�̍4{(`���C(�D�Y])�,u���<ܖkoK��������\ŭa^1�0|�o����O�8q��FƓ1]`�t*�5>ow~0�Q��e�\&)���/��)��2"��4ӂ[��C��-{:�/v�
�L�w����l�=�<yD/�ah�H�98�B�t�o��G�57�TY$�G�|p>���,;ɝo?��oi�6��8�_PD��`$FJ��t�t�.v���aB���/pe�����f<D%���MF�q����?p?s��uT�d�q��4	ŉ��>ҏs�G*��_�!?4k����?�}j�+�����G��
o�{F�PP�me�����`�G��/��I�K˙�k�X���w̽hH�Z=;z@�Ԅ���$�����FlS�����p�Mn����L4\���.���ӫG��s(��m�#�yHZa�$���Ԕ�}��PrS+%8#k����m/�
)!W.#|��}��U�����M^��e�����޻z�cm�b�r�
Dm��M�� �m�}G,��
@��N���,&��GZ6n���ۃk]&�>�l����W�`������Ī�O�\)p���,NQJus�Bcݣ�ϭ�]Oeۘ���8�aČ�3��g���)wD���7���/����}�$!�7��f(���b"�y�(�	�FȓO��V�y��*�~'���B�m�����Л��T��)�����(`���J#{��I!$;Ϣ3�!`�+Y����F��Prm\�-<�Z�A�g`��c�Ͻ��Cߧ5:AP�����K���T�o�o�|�4�y�OZ��މ ����2C4t
�~t���$���Ho���(V��h�^b�Vf��1��"���w#�����k�2J�VG,����
j�ٿ6�U;I�i����m�1�E^i���͛#�r�3�rm��al��yK�Z��Sz��pfB�5�Et5��;FP�(44|\����*������!��0�1��aPf�,Da��ʦY�&�Ь�Af��)Hq}¤���#]Ծ�gYyc�p_�v���4DAz̩�S5n��k���f�Վ������@ĩ�A�`�_L�+�`DS_A�_��f#15�\��UQ�w�l�VdQ7���+c�j�5%>C&�'y���W*�KRb�?҄�a��B�#Ҭ�.`H�vB-+Q�3�g����mqE+"�"!��H�V����ƹ��ALc`8mAݎ�1�}G[hp96��ꗎ0a������;r�C��߯K�s��^�M�q��+�X��K���Sj�	�t�����59J��Eٹ�'�Z?��<'|F7���x�&1�I
��^>"}�EH�lGj8�D��`�]���?~��ƣqQ@�1x�zBE}�󝿬��)�S1�dS2�/�ʄ�������V�g�{��7��&��R�pgꄔg`L�&�AE���Y����)�k#�S�1cE[����,����x���K��	���^v2���جD�Ɋ��L|��7n� ؗK�H�[@+��^`�)	��ےl�q�i�����ۻ�]c�J����5�g%Q�tl�zR'���!�S�/-�ad�v���:|w��,��s!z������T�tsJh���]�;�\��8���-J͘�ѹK(�|lTQ,x�ё	��1�H�Yz��%���e�qw���*#��{�\��J)M��ܳ���Q~B���8��إ5ld����j�����a���0s(�m�D����E��_ÿd����^�K�	U���H����%��!����c�ۦ��jt�B�.�h�GA9�ؖ�I~t�÷�k$�S���[�������hќ��}V7��7X�kZy��������n�!Y���A�0iPAw��dRo�RxPa#��1Δ��)�x{;�o�c�8r�fU�^P!�0p�5FD��B����q�'-#ͭ��B[ӈ0�����3y����!a�T�3��@�V�̒����8[��ჴH�V��VJ����d9���u�FYB]����qޑa�%�*=6����5�]���f5����Y��M@2�bQ�8��Ԟ�`"١<m���;v��H�JY�����p�>������8|��2�E��x��AI��S��~{�t�����"�\�W���|�ߵ�!�m��ߏ��!��������x���-��T�c���X��|v]ڽ3����}ɝI?܋k6��]2w��Q�V��%
�!�&0��=�,f}�{q%�z@٦�^^� T�<^Q��9�5�e�B:�����M�U?��(5e��:R��ӓp�>`�s�	 ��u��_�̾n��7���>����;�S-N�r���u�C�enJT�k�P˻vU��aۜT��1!֔�d�2&$U�OĚ�b�\@\q�0I�u�	��_���
���`n��T�hk�h��z�6�
`�9���K9M��ds��{ �2�ɻzG˭XS����x���J�S�bg(�n�p�U�Kر���ǈ��vt�TY�[�}��M��On{Zo�?��}0�����7�8�����;�/m$�"��3f�NA���B���wP�QU��kȍf1�6��#G{ĳfW8��ׂ&�A�Z��f;N�Xe(�p\bg��6���]�5뽖��CQy��Y����ƍ#ԖP����2J}C㴗y��f���5j!��r�|'@Rț����V�e 9��,M�T�`n`���?��c�h��H�e��&�9ZG/ԙZ�a���:?�M)�N�Ȗ 4�P	cu_=��w F$XnT~L�>A��}B���fb��L�8u��x�߻�tlҮ�%����
�q ��4�#�&!�+"n�+������҉�
r�x-���z�w�ga�b�5�w�^J��(�K]Oh�]��efco,�8�`$���h�R���4��� '���{�iS��5�0%������ΪY��B��Fp�o�n�W\���(�se$h���~v�b���䜌Z�:�{0��>�(d�G��J�=��l��0,���r�R�����o%bB(x�1�� l������"�f���:����zl���*H�F��\�bO��%g���f���1�WV4T>�*_���S֤���K����|x�G��i���m�J�m���^,���w��=������v�Q)F�ɤE�&x~]�I�>o���]�T�'	�5��`Sv`>�oՂ�����G@�Y .1�p������b�A�	�0?�0h\��c�c_慘9�r_�A�m��K����Ǚ���o��:�m|T�9m�[H$��y��@)��Q���-<Z��?�ya=����V��5p�%M�4s���e���qTM���?�\��v6���	�\�����ILD��ʮ�\���g����/̤��_-G��FA][_:�31hW�G0�� ���S�\��ڸ�A΍�8��W;���)?@�5����}>�`l�-Sp������� 2�"�	3����%�`���e�`lŹ�7�M�#T��}V���1ĤT��"��H
C�uϧ~
���A�a�A`�q�uM���c}��7���\�1�%YOX$	�3��EŧDa׾��aA]^� 7JV�s���hXI���.���9늬�N	ʻ#o>\�L��i��q��G}҇G�Fys�[�lJv�<)��F�d�� ��+ܵS=�'õ�rͤ��-V�� ��)I�O��6�CɏlуE}�����=��6qP1�#oz,=��y�b��y]Ƀ�D|��f�|A3\n%6�4���9KաӀײ�޹�X�d�L츋������- ���Ɲ�[��{ւ=�Iv4F�&<���7= N/^��{� ���Y���&�?���"��Y�zF������j*�tJoqQ�N#zǉ<U���������4�[��t�p�!Ic@a//}� <�"��������zV��2�����W+S�(1�z!��'2[��d�YFb46�m�;���$�iA�Cֿ����e�@�u"���=8���"���]�� 9P��bg,zמ,W�^�,6C��x���QX�i������}��"��n$�&[��`z�NH�e,��D��Ym��mx'i>քbh٠��`CI��6l
α���LGq�zE�v'�ݿc��o�� ��\y��L�=�8�n~ND�z�P!�[,�a�����2��׉�e@ZF�%���ȁ0�~g�v=�������y��ڗ<��r�Z��a}nLڛq�V�)��YVb�)W�.��MXلX�pؙ�)m����K7��h7თ��q�Nq�P�ٙ�f�����`���a_��^�.@|G͚�R�`v�9U-/K�n�f�����:f�شJ9(�.O���ki>D���W��ck?�����6� 3c몸�����p {ޥ�l"�[�;}�/V�P��^���8���F\��f��"�Զ3u���*XL��9�ʞ��7��JR=y��9`���J���)� =��RZp���_��ݏ[�
w�3h�P�dԗ��R����V�q(u(��3�o�0�������]�zE�S��4�s�R.�����g�]�Aezv����+}u�w���N�r����ϟ�a8�=�\R�s\�G��!��ʜ�8!�-X��S� �퐲<����(�f-\#�a��U�a�a���h]�q �88[2��O�E�����U��ROG�6��Kg��?t�B��� ?,N��6�ژq\.}������xM�����F�T��wz�~��e"u_�D�犡z���9޻�؉o8	�x�3��悈$D�a� B!��f�z�X!3'�]��}�*m�d�!+��G=��R�	sru�n4�{z�!qy1��������C6�*��0����?-jS����}84�B^�<c{[�\$�;p��X���щ�<����π�
�����sTnY27"������(��Ob���kқ&UKB]:L�tŇ�H΁I} ��I��K�,c�����o���!�1$�>h1)FL
�~G3o��e�M9�&_5���*hE>d+�"��Ċ�D���l�Fǜ��#�e8Dl6LJ�|�?�&����R!tN��	�n����whp9{���S�n��R��0�/�{ }�����bYb�c6��� ŗ_#�Q��燎�*z "h��) �'0���Ľ���y���D�a����'���[J6��r���߰��mKG��-�$��?�=k 6m�ԃ�
!�5*��`����Wh��ݿ���d�����xzd6F* �l!��#���_�ٍ�y����x�L��"%�vo�̶n��YGJ��^�5&N�<t
y�m$	�&84u�<�Q�9('5��%�9."��3���D�ߠ)ͤ@��X����2n':&���h*?e�Y�zgy>���.5�F^}��	�"� ���F.�P�O{~i��^�O�fr��x\�&p��g�M�pj� �r��Y+O�Fc��q�\�hq�T�9x�B��;�4��}�"OO0����c�J�A����]�&�	X������q9�F��n�u-�ݧ�F�"=����#��kf|X����V��6:s��ӧy#',��d}!�.�8����+�z�S����n��6�����S/½��gN����#d��r��8y���?��f�CZ8��j���\Cp�lI|rA3�\�	�Y| ���$�;D�>�پ��U�|.�wsҭ��"U,?��	��--�R�

p�k����O���:yҟ1�q�c9��S�KJ�X��B��`MP�,����ok���Z�~�C�v ;��P{Eϛ���� -Hv��cR`N��Ne\��'��<_!�]��1��c��a<�g���\KRy�t�+N<�NE����e��WB��X��3�� V�@@A��X�c���@�1�WY���i
��e�a��?� P�3L
y��x:��0Řq@�_ĸ��*:�2?���"�U�k{I��kb���u$��R�QY��(��I�H������R)�;����,�G�kkɮ��ñ�!L���4�-^z�]��7+?�+��om>�"��1��j��?�iu�3d�2��캿6$^P����a�R_��m	�ƛZ7�+5a�P\o~ѯ�r���oΣ�QyD�G�&D�N�x?�DGc��[EԒ�F���_8뉖�_0� =
����윚����^�3��)Ni��6 &8D���K(u@6�O������uT8[���<ذHF-�~u���#K�X�Qq�� �>�P��#�f���G���@�i��+����J<�Gfp��\�+�0K������3Q$/�R��W�:#r��ti�ʃ��!�^;xh�܏��8^��M�aR�CӮ��#���uU������W�ۏr�����?�[ɢ�$>c��U�P���Y���ð�=9;g}V��j31S���6���έQ��6P���̸	N<G��%���k��+L��v��(3tǞ ��k|m^�6r��D1r�hC_��^��+]�%d�S��	�P:F��	X��I�'�@���������oП���Y�&c(�*��yUm0�	O�g�a�.)��%�(�晃������%.�߱f�M�(�# \�<ӫ�`�	e��m�E.��\6d�A�%�$�\��9&?�K��c*K��6 @�`�y���Nu� ,��,�\�
�k�ڬXp"�Ӂ	J����� د�"E���h].^�hA�:��&-��&�o��z�F�R7,��9�]�����m�C]��(sN�i� W{�Q#T�~��d]�+
P��Ĩ,(5D|s,w�֗.vS�:�m���/uI��i��S$�!)�%K~)�i�u9�Z�p�o|�G��D���e�XBo�~�����]-�P��~��k��[�rk���dU�	I���	@H����6���Hw7i�yE��̻��2ׇ�X���=D^�2=��enqETM!��/8���(C�g������_��@�����v>'��!�P�R���~�r�LRΠ���sm��a?Σ�c����w�Ȁ��>yu%�z�JdϘ���/���qE���p�,?�T�L�"R2�-��� K� d��Ա�	�)-���!zg�Y�©D&���
�G�Z<|$�.�����Z�Z���I�T{&7�:�
�:I8+ '�Hu�7�S'��J�dVƕu�����a��k4�V�����B��q��(���}��#9��I����F��=�F�)&D�^�c���\ƅ=d����Bh����j	<��4��ʛ w�n���f,��u� �"�&tٿU�����X.�B��P�nn;(�M@��H�m�l�*����%/kn^$�� Ԍ�K�Z5N��N���0��v��ji�n!�2<W���k���X�Hք ~�>�Fa�Ǧ�i��fRx\��@ʙ-<g�j�j�|�	��J�D�0j�lڻv�v����h$�xH�����'�PB��ݚ��<���dwċ<b���9h�Wd�JB"`��U�reL�Ԃ]o���[d�V�:q}�م��X���az�e�a�[h�o3������Oy��5�<��x�6��V�����?x�sz���a�C(B�� 2)������'��߾T>� �yVV�ڵ�f�B����n�=�D��l5  ���H�dZ��)����h֖-(�����W��ܳ���<�6�{7A^>��d�۬ҽRhP��2I��ɟX^#=�_����](ςR����Ux�-|�0��EXA�"K�:�A�h�~��P��{]z�ڱ��2lK��>z�˅���$���D�ԇ��T�\ኄkްkE�����ٽ_I���Z�\�{�	�?����/����OBBD��n�ܗ��?���eY;U�/r?[��5$~�B�-5��|��J����$�f~��$�u��Pu�x:� ��҉��nI��_�?�8z�<;>r��9�I�^�9Z�AJ��[��q�n!=X�nJ 720T��چ� ���y��cj�-Þ�9[�yh�a��r3f���t��RIc~Ur�a�k�����Q!JfU�ŵk7�����.U.�#���m�+��u愬������U$����w�闆ɀ��z���N�ʘ���⨼5�Vb�YY�%Khp8�'<�}�v�,O�M?i�l��]�����?���np8�)t�����5!�M�HS�j4b+���+0=x+��*zءG�o��2��o9�T����S���o��^t�7�#|IX�G��?�TbVG��5�i��HT�	��C7�!�Ga;1��a9��|E��I*&P �]DW��0µ=~^z�c�#F85�m��-e��i�y>��Q�m�U�Dr���!(���x&BR��TzA���w*؀OŁ���6Ơ���@�\�G�.�'�JgjM��f�l���i���,�é$� ]B&��)����E��g??N�#n��P���W<�`�Q6Y�����Ѿz1��D|"�fd�x5B�J�.}au�����<�R@��Ƭ��
�ꗐ��:)a Ӊ��EI�^�)<I\1�;%�8�i�� a�b��L�HN�:��St�hSL���6��7{Z
ݞ9��B��]��ȸ/oH��� =��mu$�F�)\�*��D�g����U�hT�
��ru��F�MS�\�m羟"D�}w�}��cRZ���/u[]���c֮}������E{	f�u�|���?��+wM�jm�!�b9,�z���,�����/8E��?L{�Z��s���sB��z�d%��[���	$|q=���6`	�y�����rh�����JV���}}h*\ ���W/�!̽��ԡ�����I/j��J*�o�������8��]:�����u-P��Z�S�o�D,��B�f�C7����!KM�&0�9E�^@v}54�9�oЁy����I#�/+�wzJ��2��D�$B��H�z^odW�r�4�QץQ^��p��i ��|Ua���|K@7Ď�&��"� �z�tT* {��K��o��J�<�X�CF�{	7�š<'j�>,�(��d$HC4����[>ќ`u������]E�
��%+Q͜�b�َ�a�&k'�$�����m(���$O�}N`pF��g���̫�X��<X�ra�Zs���	9_?"�gO]'@�����o}A�u���K����U,�8x����h�-��㨊�L�@�&�k��S�A?�eQ_"Hږ�t�G���>�����G����[T-DEg֣x�S����xz�U�|0��	�1T�X�+�h�
�oCB ����l����ɴ
� ����N�]}��	�������jEL(X�"��"���}y�Y�D�ó	��_�Q�H�٘��}�봼�q
R��)G���-�p����8MC����4b1+Уr�'#-�k 
̪,d��2��b��j?_���Hm1F�1<�d`�{�HA���.�����۩���V��A�̽�zY�ꋞ��Q^2���:�|�ܮ�	�ȯ(F�.>1G�G� ў�~�?�昈sΏc �K5���'&��<��}Q=i�����k��Es�d��z����6����|��'@�m�]L�}��7�xx�]�l���ܹ�ro���7⡻l��ES���&]�AD��P��4ULս��.�^�c9��67!d�6��y�J&䀱���1A�����T�O�= �*0��-�Ҏ��m�czalJ�:=�$ec�ʣ�-dF���3�I�O��Q���������2�2�3<�"�=}�!�
!E��x����:��ڨ+�R
�į))=T��Y�G�;K��[�«��fn�I�Y�c�y�I��0a���j�H�R���^��Vun8��!���^/	'��3�E����-Nƭв���O�N��~1�iM0H�������/5`q���Pi
�	W$y��T�`<L���[�W���"�K_��F\���3�cr��rO��a����'
\��q�q�M�k�����f����8h�s�ANM�)�)�j���l�uXA�~���1aU��O�ޔ	⿁0W���f�3&�������E]���h�JW��������=2[��H\z?	����r��;vk�[�n��F=V#��NM���iu~te��f An�^��Y �a7��;Y�,�v
�n��3`jN4�#W�Ix�}�+�{��ԗ�&�9O(�fx�v\l�U��������z^�7_��F`�,L������tg����~h�A�ME(H�	>������Lb��,SJ�3ਣ������_.O=ә4��ٺ܁��r��i�ٝ2z�keY���&椟� rX(C�*z5� �{_�W��g�/L���P^d�h�;˩�bp�䛮���P�"��?������T2�u��t���1E:�ѿ̠�	��}.h���I�(W=�&w'���ԋ���G���G��lLP���ʉ�Z"�PNﲤx��A|v���ܪ��	7��,����o,��Jz��{P��13���[�������Q���i�pΞB���oh�'�:������g �'\f8���,�MJ��Ƅ���u��zu528]�<j3�[���>��Ŋ��31U]}}���������ˤ��ު4|*/�͟޹}�ڭ�Rwj�M"�Yv}�QJAYa��%�nj0瘅sͨ�P y\
k��lW&�"��Q`@Te/6w��"7HU� I"ɘ�����:���3&�K��ӂ�����Tܣ�wԐ_�5�LRo�j�~����m����F2s�B�B��S�����cq��A�D�z�1
=T�K�@��'U#P����I�^�x���f��	=�%&��á���;r��W���EOhNWJ�n�ߞ�)!�	q�qF�!@^`��B��б��/��{��_T�G}4h�И>']C�L�����A�*�XW��=���TGSsN�>�肯!��"�΋L?ķ����L�����=��@�3J���'1�0�g��#5N�J�A��z��_����7�З�?��?�i�*G���)�ic�'�^Y�$à�C�������#���0��ޒEv@�(�5|E��9���l@�չw9,� ��uw5�A�������Hm����8��ϱ2+�������N~�p������A�hnB�g��w� ��>�V%`��ۮ�9[��i�q�>؃"���DuC�+7PAU�:��ex}����ZW1��5�/�j��������tvx�ߑ4����ؘ-�� HB��M���=E��dA�0yc*E��領��[��:kt�� B,�C�?ޚ ���*N[�n��"�9�����n;�98�"q���kB6D׫���	��h��F�		sFIt$�03�,��>�A��D�;��Q�Z�� �B�"}�g����P��I�,� ^T�ʡ���uv�����C��7����R�'���#{�mȠ�E��+�ǂF�~I�,ۤ��> ��9I�#�ǧ�i~�(�L�ȥ�*<�4V�2�P������(dd���--�Wm�|��פ��vPŌي�,�>�*��O>�!3	d
�tRȿ4��j�Mh�h\��=]k�K����]䅥��̞�7��3�j�зŨ5���t���5Q/ݱ�+����R�EAWO����~�a������b��-rmYq����v�H+����]�]~ݰ��矔���"*�s�W��9g��[�"�x���)���2�m�[5��.Au�������mKA�����#��:D(U�0r!�����k�07��Ա�����vm�˙�|5��X{��и�i�}	��]ªx����'�7��Կ���l@�'��a�+��8[�j��2�&{��
�>�tkA���t�d0#�zb:<�!���"S�$a;�ބ��j�4!���{A^6y��!���4iև���7x���Y��($Ék�z\"Y9��K<eX�GK��@�8�cUr�yh�犳XQ�����n���"��I}�е�a\��87�%�X�̗s���}��6*@������ʹ������Z#�b������؜��zF~�䏼D���pXIYD���h�@m���>F��҂-�%���6fl�ަƦq(mt!A��3���>�����v��!�)�
���@�'��� ��i5a�����l�ɂ�\z؊ss������ڝ�}�o��X7!b-�B
��N�=ݘ~��2�]��>=�Y�����SB�����)��w�4u���sl:���Z�F��	t����G�c;�3��o��x��&��E�7�kQu�����|��4��sM��	�)�~z�_ڌhV�P�{>hDo�ث��wT/��\o��.����P!$�7�g�y1�D����P3�}M�Si�_��ΙU��@]v�7� �t�0�\g��}ش�z��������؍C8�y�K�� �A}�*ؒx�bm�7�[��u�i�`H��r+�����������#�B��W7BcG�����<~G[Y�i�Q��A&Z�m8JZ����K��~��W��V�mҽ,��f���*ؓ�S�P�ڳ��c�����lɸ�v��<�>��_�9ByO ĹW�5�X)��):�Qd���Q��]���V�w�	���G ����o �f��r�E#!�������[}�5)��z4L4V���,>i��@\�:�8o>7-H٘�����!"�h����f���?�|��Y�m=��>� #y�1��iQ����E�(��u��$���v@�'#.5k�4���N������0��x�7:�!C6�����U�'���(,y��4#@��&���y�`ذ�n�������������,j(w��a�B��5�r�0�JX���A�8q�v;�2ȏ|�Ͼ�TMJU��vj�s�И��I<1��B6+�a�L<U�&l��\�hkA���4��s^;�A����c�U6W�3y.�u���%n�H�0:lm����Z.��)r�&�o?D߉�9�V�=�`GkQ�1ݓÝ��#fN�Lׅ.�2~mi��`1PO�,Y��ʛb��5(�m��rD�̄S7��".$wY[��b��-UL��˨iga1�cM(?	�_}ޚ�!�e�I7���L�w���#�i�R�t�"��'��~�3>��@����=�Z\\�E��',�8S�,��\���^�C����;�iJ�:k�z��I!f��E���c�-w7�I
�I�����%}�ӧG��D���+>r�Ɗ�+�_�>+�e4Pwk���r���xmF������՝����m�*��F5��$io,<�+�'jE{n�l����!߳��{7@���藀f�T
ź�²`k"��w.�H% V;��;�~~%0C��:�Slχ���9�C���s����]H��6m�Y��=)V�E�����)�<ч���z�[{���~%Hl�db$�t��A�[	�Y�=8��7�CV�<����Wd�?tҠ��}{{��E��_�l��6,�Q52�#����@[���V�f랡7>���#�q�:��Y�����]�˔H�@>�a��o$X;'@�[��sF�P���/3n�lo:;�-��B���C��oFq�o��ۛS%�<�E�Np���hjlKX"Y�z�jt4�#�۪�'���G >����אf�����1k��~&�33�;s��3��A�]�P�/�o����W;��s@��E!ӒbO{�W�S�܂���>�҄1{��|�5ڴ�R���*�]G�B��(G�����+�������D9���1�ہ�=硈 �i͘9�ر5�չ�o�$����S������7�R�L��~��I���	j�-�l��N��������zM��]����q,�G�XcpGlOqJ��h�eEZ��� ~�{��jԧ&�cTK��C�]��m(�q����l��%�~��;������Y.M�dښ�?�M��>����`$�K`y�%�z�7e�\�r��e�R�;ڌ:q�����Ie?��U �Z��5ٛ���3c�L�U�#�r��Z""k<�ޡg6_���>��s��k��~�&F����L���Yu�	����׊�ӻ�� ��֓DzW�g��a���ŋ�c�@�[�s-$�䰩��N��~�?�<��%�����yw�����<��f��{d����H׉�����/}�>Ml��؉$��<���ⶴjp{>�2ײ
���R�r�����uZ���u_���"�mX�d��U����fۭ���,�O��6��@ν؋C���%Q�J�]ڼS���.+�EydD�k���$���jT(�MOl�6��g�N'�E�W��T����)Gw�2VR�BXL�^z��4����r\�����Ͳf�H[��A]4^R�v�''�l�b�e>]T��p��{���p�/�p�ah�_��e�݂4�Β�_�sod(5J�T���-2y��!����� �d�AY��6k5�aw��D���WA��"H���^s��ʝ���> �$�m/;I�w�~T�YQ��S.���^V�|ˤvGY�Cb���#�՚�8S�4�OLA�c����|�48����D�T�OL�d$�4�E��ƴq��l.���eT��N���p�������wW��:[X�	�����\[�1�Z�s! P�m�����2�EU����	`n}k�xT71���s}8c��*��>������Sbs�I�H��#����u�w�ҡ�+��9m�`)��=)�W�0a�)�$eU�#����X�}�Ru��:��@�3_�m�dH+�C�G5�?
��1jۈj���d��0S^�%L���N��'�6����Q5p����<��H��`i��~��Ԧ^�Aԛy+b�A�˄Zu��_��AF����腹��?��2�'�è�x!k1�+��'΁)����eY�X���k�BW���7�z�ʌ9�����1�X����-�F�����"�۲��Z}�����l����4�y�Hsx"e���W��[��N}�d4!k!�tw�?�n��o9����Fz���\h�4u~������>�:O�l)��^��g7���K�DuX�@/~1W�}4A��xL���8:�5��T�n�g ��_k6�}pH�K�g5����l�:�����P�<	"���Y�����n�Aj7+v��HG��;o�\��T;�J	n�@�͢l��~��kj���� ᄴ�o䐯��	�@�e����rX�A{�≱��U,�zE�8`
�H��->pI�8fLQ�h�I��嚍#ҭߠ�k"Ι2����lX�$�}��4������g0U~;N�Lk)�<b��W�׼����a4�Eŗ��It �r-/{xC�6������:NɅ�0�>N�:>u�E�Oˁ��m����v� D^�"�X�@-�J؎Q:"����.�u+C%Pjk,�h���Z��w}6�wf�b��k�)�$_��q���.�]�<ʭ�:X��j�+�q)W���ݲ>��z9-������C�8��c$�8��°\=�<���H�o�OTqAе
5�~q��m���>?o
�1��j)�j�����Oi�'�}A�@j����"&Ӭސ�s�t�
���Ӕ<L�C����.��G�s�	��|��I{���J���^⷇ަM߅���l���Qxգ����
��  �������O_ԌB�����d�Z�����}J�7�����]�9<�U$6	�p�Y����C8yXQg��f32�Ju�{��d���7�_�rFQ���+�߆Dɠ:�4�/=މ�6g�*�j�)�u�
��臠ꀲJ_��a�w�`L7o�U��.��?��W�W��97���^��B���;�ϺM�q���'j{�Fo�偸���c��Wv�j|��R�ǖ�8��ދГ�&W���	�7�U��E��,���@�#(��W?��N�Z�S��_�U��&�G8�0Q��Q�0 ;*�vPY��9p^�C�p���a��GsJv�C����]�u�[��~�̳O�4���MY�-�+gBX��4�vLHOq�y�K�����'���%�Ӧ��8��w�S�]WZ��zk.�9�8!�������s�~:f�<��v��/77s?��J���4�}�����1��cr�0T�������lc-p�
��Bwc�>�rX[:���6�4�|��q�7���%�w�*s�jM8�g�����{0�e�5��2 ����kR��B-�E	(�!��opv��%��d���y�D(��,�)�[��Mn?X&(�$0b�8�ee`%��$��v���X<� ��%5>��R@��z�,�O<b����˜��hR��=�>�<d���``�iMzW�\��V����'�F?b�v�Ж��"Z햞G��~6~D��#!U�Y�ʹ������6�"�q�(^B��{Ek��+l���a���Xa�v5���<���0Z>�}$���;��E#{�*���A�p�P��ό�˗�����R2q|�ۈ�Bg��h�����+zJ�AS���z@o��g5:�ԕUM#^��۪�����������j78�we�� ���T� J��-zFQ����K�
E��R
����Fq�)�a�wL3����!5>Ԅ��K��%8�):�yvT��*��볃r������J
K���w �� �RN��Jj�
�]�N0 ��s��
q����g�	r�����:�N���@�%0�^׺��=���Q(�ӭكo�F l��lGD�6�����b���N)�Ы9�:�͋}�[����7�D�K����I�{����%�i&�=�^���iO�v�CM�)��r�浮CCNd��w��	�4��a�|�^"B�.�2x����zv�e�:{AZ��=Q��vlڻ�3?�0��MLx@�7�J)���ݤ�����'ꢜ��b��מaO:䯞�#�I�r�g��h�������k�>1����9i�A���$Y�T�O�@)0� c�o�$<[Q
�pRv����P�J���8�g`ϰ�ȵ����ـ�ƾgм ��������d�����/�D��W��D��5,2�QZ�vx�]�c�ҹ�ix((�O�����\������̵Y�笑M�R��`Q#�
�I�h�n�M_�tA��R'XmDE|uS&������C~�C�ܟ��_	�Jg��%3z7$Rp��KEx{x��,�-K���������BıE��Q�5�t���������u��E	`ᰪQ�.����+�|�J-�Y���`#��v%���R`����s��F�^�9�z�u��\ܩE/Ц+��DꞞ��D��o�a~��*�$�kv-��}��6wm"eDܘ�[��D�����E�w]�I<��=%yⲏ�3r�t��N�I�K�k��N,��VZ����C\�٩\�Ad3���V$`1{*�8��O��B��F* 4y����#׈�]��FCdn��2��'5�א�2���S���Ճ�u�����'C��^ۡajC�r2e�ܸ��k�C�b%��UYT��<���^b�ʓA�fc�^���9XbMҹ�i\��/>��߾A��F���(�wN���0�a֟�~d-���R�x8�Y�E�dP�vо�h1�/�����nu}�x2y���;-�e����l�N��J�d��b|�l|=���4�	��+Y7�:n8
����ܗ�o��e/��b�f��y��jI������]l��L��}�}p���<}>+=늱�� ��үK��+P�t<��:��ܰI&�4]��p�_.�J���X߽�>aGv��I��w�F+Y�X�A~��"����p�1Z�;�����etHu
H"X��ǋ�6�}?)O������Rh%�^�R�+bJ`*�\��"�����O4�����Z�S7�bA�
b3Gy��r�/!�¨�~�$v�G]����[s ��k\��z�>�����U>�܅ڞHr\�F05Ɵ��'�������)�m��l��Hx%W���/O��_K��f�63�DJuءP�|-�,�=�Jg��V;���:ܮh�����Mw���������c�A�pb���D�/���ȸ���{�(�?pCZ������8�<~�[�Y@��V�mG鎧R8DMKJ��i]������`����b
�M�}"�V��Ll�b�11X�/�Ez ըT�Z�NC�C#�֤�3.�*;a0B�B
� �킉oۊ-䘧h��>���E	j�kr��9�kN��S��#�� ��*�{��K�N�v��w1` :G���+�L.��[q5�Fs�����X\�=i����CriÅ��_�I��2~ri~�a�q*�@��8�I 5]|TFjK���A�g5����%����_?Q���<��Y6�0��pp,v�ѿ�ru�Y����E뷓	�R��b�e��L>��n����b�
��<�9;��B�o�m���3$)��4�'��~Z\,�������rn���J|
L�������s��%9Y)�!��Q�^�Ce�P�@�߁�J�����d&H�Ɯ5�I��NFp�i�����@[���\SFh�H�]�e��T���Z��f���C}����G�9�F��^d;�DW���SE@��?d�d�^]�GE;u[��y��J�o���f�o;�ç(%��]����:Wܬ�QJxe�g�P���h���
�����
�˙�tIK��R��95��[-�aי�*���r�/ɪ}�8�Dܸ�ɷ�"�u��y#��-[D:�_,���ٜ^V�.%���>(`<�zPS/&$���F�����Yr�&�,Lx��S�{*�n�?S��kcfrw��h����Z�)	�['P(�u�BR�Qh�U_箨�Q S폡p3��f����y� ��	��~�?3�KS�M]7�� ;�ayA�CTf�	r�;��"�!'K��tD�0[�x`�?.�f�F5bꛭGJ��]J�[հV����|�:�����'fØ�؀�������&Qz	|G&_'$���0�q��鞕dP�ǲz���#m��Z�ș֢��kC�N���jJx�@� ��#�	ML��I����P��:c��m�M�ۅFG��"FsG�HG�G���N4���u�ߏ�KmT��������C0k�]$6�#�9�u��ʜ�
a�'�vx2)}[��k��à��<X%Fwz��)�dz�my��Ml�iV�kۤW���Զ`����*�5� ��D�#I�]Y�/�q���2�_<W�im"�y^?���.sYkkᛠJ���na'@L�������b��Ik�������P� +1f�*FL-a�ֹ��A\F�-K�%�����=v�"1�������/b�-s�p��ٳ�>��G���Z�Q�dY�w���|���fS~�lC����4�h> ]7.FBf�{�(��1$@J����_�3�E� )�����d�����oY�3�oш�i��5���d��#���^�	�Ɛ	���̔Pe��!�킵	���q�fk�$W��@����̓��I����۽�Bݘ�v)��
Y�x����t"���i]�k.��ٸ�b�(���$�SI�����.L'�~!��*.%G��h�?�vݏ�8��	��퇞������V��Zż��[f��|
ߊ 1`�X{�+}��5.σ���F��A���c�^�qxG��[���W������#n~�	o+IXG�q�°�x�̵��Z��[�4�9i� )3��k�{�p��\ŉ'�4��������1g��&�!;>��<�%3�G�N���}��ս�0�7 �t�BG��K$��7�'�/3|�>6�)r�ϸCE	�K
�	�H!�慧�x�w"�Z���-s`�c���o�Xٴ��B����"<���kb�lxr�I
U�Ed��G��Ŵ�LP�^��������d���``�7;^��ܜ	��_(?��E�����U-4<��I��A��lSiط{)}x�g�����R���T����n���T�:���B���QQCm�j���F�ֶ0W��Ȧ��╅��WdT１&�u�y�.-I`~+15��b��/��뗴����9�����>c�<Cڡ2aCN �� �J�0s���A�x��](c;R��a4�9�'R�\B3a�Ė}'����L�u����ACh�r���0�Jhz�	�����\�e��i��Z�x���̯
m�ߟ:|����>���$V�l2�16S���A8��SJ^'�D����}��s惈U��O�՚��A��>K��R�P��e�6t�4���b���"��Q�C�LC��Y��D�f�-�Q�����Γ`�C6&5�T�m�E1H����@p~��э�����`�(�d�bdw8��g�%R�g�c���\���cI��'��[M0P��=mCH�� ��l�v�+��_�E�g�0ڏ�}�˓Y��g�W���L��~����UK �ԗ-䳍�W���S~ֲB�����
�S���豊�V40�Ofl�T�d.��MC-�Hg�b�b��&'@=P��گ4.���iR���b0���]t(�wS�|�f��%��o����K��, ������g@����lE��8p,�O��'�pT�A��Z�h6�[�>A*�"=}�.ϟy��-D�,5 LGO��h��g�����Z�tT�����:tl������Tuh�W�O�^�p6A����2&��,���D�2�U����KK_)ek~������gN�KX�<]���C�}�M=R�@���I�(~�%|��g�������v��H)��Sw�5�S�&wN<4�����R/�.gŀ�����{�*D�rR��aH'p�V��I���N﫠���Bٙ�ŧ	�'��y|y%!~f�۷}I���*�e�?�PB���L	���ܷ}ӥ���=���{:1����r�_����ɴ��b�)l�M��8�0�c2��_��G���D��mX���Q�W�H�LT������8�D�*�#�ME^��ѽ){Vd`��Z|��jPp��j�$N2u���$�"�A����v�Ԗ�9@�߳�+�ԅN�55~�X��W�U�@J���<��2��&p�"�3H7:B4�ĳ"{+�җ � !޻-6IS��60`^���RH)oXcz���������-CG>�.)w��������{Ė�y:�e���{Z�E'\H��#�O|5�s{F���ֽ��d�# [`z�Λ�<�K��Z�7�x��7��1@��6W�?�mKD������G����y�>/��a�/����R��A��;�\���$���<<,�\){сZ8/g�K"5��?��-[Ǯ/�,�U��@�
 E� �)��JK��ܘ��n�D�'��۵�p-�v�?��>��LΫ.��Jd�U���|l�r�z[@�dC�Ϣ��h�\��!8V��^i��%�TF�.����%�朗 v@={"=�ɩ<=Q� ��7�"���/v��)O䈭w�h(�q'Z8���xB@,F;	�Бn�T��#V4ԫE �b���	�o��L��2*�Def�^tY��B��a�T ;5P�5y?G�	h�Wt�K��q��:C���L���ѩ�;3�p~闏7��_�"�����znv���m4�r+�&L�b�}�d@/�"���a�R�����������6P")���64��O��
��Rv��s��
S�&g��>�!P�V	lj$S��0����Z_�̓k9a���*2��U��!��`���~^pgI�Ȥ���$*ƭU>����k�AP�.�E�#��_�KS����1,)����_�X{U�b|R��������0�z�Y���
ʀ�Z���7;1�!��aW�IQ���C�8���;s+q��Ѓ@��끲 O5��4�����,���`�Oܳk����f��u~r�T��R�du�F\��*�s��˖�+��P}�v��'��wF��0B��"�.s(VnU���?��	�iY\*��R�꺃�,�o�KZAn|�b(M'����T�ׯ+�t#���=��a�P��QP��YYsο��$�><#wY'F��l�3�2���俤/�U�2r�sQ������!(S^"���[cꠅ@�2�aV�L��L�i��w��ä���Um���u���m�a�UFk�j�s�0���Kp�n'�g)O���6�8� $T�ɌCmJ��r�CX8�}D�$�^�ΒƠ��"+�/
ӌ��D ��?b�bv{iH���;^<�|Ђ� �xA�Z�D�o���f+�vA4�҈�PP�ʒV:2���-2υ�C6V�e/G���<st�{�'�jXr1�#S�S�f�	��O���rxU�=��m'���os.z$/�0�d7��zb��}0��?G����)�:�y��t�����?�7�x��2S�|��Ǐl��/D5$&ԭ��I�d��p��l�>KL��?)XRO|m��¯ҿ+�1�j1��W���0��'�T L���T|WU0_�.�D����`���Q9�-��Rͮ�m��V�)��g��q���h�(���d�>�d=�9I3��\�� x��j������/W<�$��N���h�1�E,2�4�P?�[B���u��@�**��x4���t˘�
=J]�k�M�`��e|��I?��Dx.py��#�G?y7ima/�u�Wy3�S\+i�2�������揂P��)
���]M����ǫ>2���\u����ޛFT?�z���S�1��~S�\<N����B������~蕟h7,��!��Z�d��JS�~8����D�u�Z�KC��8i�	�9���l��i��7.���h�h.utw��M쨥�J�g�<�
g���Ge�!�ןf�n"!��HD��0,�\���ጛG̺"�Z$�#�u��^��K��Pk��?��g4�_�S���*f���Z<hj m�)�EeZ��u�ۿ遷\�ܱ��F[Z"�"Z��U��(t|���H�%I�����P��Iq��!7�6�U���~����{v��p/0]�����,��8� p�F���T����(-H�N���II�J=��;yƓ����4.p��
���2/M q@��m&\�|����{L�hQF�v���Gm#�ne���U� e��flI|g�����6�G�n����Q�2n_Pȃ)A��N�-mCd�����B�����E�����t��/0h�UكQlvW&J�r�����8K���,_BQ����\Ɯ�D/Ò��>Ӂ���A
Eک���[�`� �5��.?=�C��b_�9��6�J��U��z��:���J��_n��A��f�{��$��Y��vxb@�'���V��J��{0�W��J0�z�����v��`��D0s�>-�bo�O��������4<o���]�5�s\A3;�֑��4� ��oG����A9=* 9X��xel:=�0@��B�����Wp�O{������A�m����!���Ϛ�U�D^ �rO�ށ���W�R�n�|�z*X�ewO�vˬS�C�v��Q���e��o�p���'yd(��z3�6#
a������S�u�&׺�}�)���H
�T����*aa�Kn��W�e'��S��U��������e^���wZ�8�p��8���*>�����> �s�T=sH��?�[t`TUWhfJT���l����vC��͠:ѳBV6�iV}Q#t�k)���þ�[��ʷ��y�o��a�����ǵ�*d.�q������k�^��=O��� �� ����5��CsOc;�+p�BH�z�S�:ᷲ�����El'�~m_�L�` 9�r��<\r�s %� ��3�~�V�Ъi���"��(v�g��O��"��W�D���`�*��ؐ�_�-b��ר\��٠o��ꕰ��;��p)߸�ćq��,n�_�ޓ�A�7�#�mܪ��x�,�HX �x�0�L�\ 	"�����k�T��)�Qų���'��GG���ƿ��-]�Ċ�p��_�~cc��
��ͦt{y��g����O�~�����"�wq�
�aj��H���'+��l��"HX}W�T.��K�y���= �`��Z)s���C��GgO+A��7���G=�HR��F.�(�[cn	 z���|T�dIFG��E�D+^�����|��Yq]��>�(i���]c���ϔ��je�֘�y�0������$U<��a%me����l
'�8Ӗ��_��V��WL���Cb	��x���[�3 ����>�R$u��5f��("��Ď�zSz�X��w��744�֠/i��=@�e��"6'��mF\���:�c��~���W0)��0�$�^Ŵ�p�Կ9�/s#�"o��Z;'H*���+'0����.Qj���n�P����⠾�1����D��Y�Y��� ~\xfg��ɞ�v��}l�a���G�pDbu�oQ�5-�x-�]r�ȃ�0��G��XǺ�2�}�(v���G���o����\M" �������Z�b׮t���B�-���j�!�,�x"j�H�h̀��A�yf�e W+39Hf�I8��0ɦ� �$|�5h^l&p_���=���̕،?�x�g�6 f�[?Ҿ^q�oڧ�8X��z9�0Q����/���J����3"L0t��t�"���/�PhiH��2�H��zZ� ��J�b���W��F������N�k�h�`�a�����+I�m3���=�O��Vs;)jr�NE��Q�v�x�$�!=��[~�}����պT��>x���*�Q9�N���ʭ�JuY������w�h������ �8��rIp��+�b���#�SqI��{K�l�.�j�1����׉,����	�,)�)BnR[L$�^?]����<Sy�Y�H� �8q�86�W�ufF/+��}Ӿ��P����fcP����-21���;�w���X0:���n�Rd��VU�c��^[�6��z��`h��G�=ҕ�s�ЅJCHP�Z��:����ԧ$ڒneņt�aq��х o�~F��u�uK����5|�C�Ϗ*�_(��t4^m�&###=�P}��������'�q�u��sz�P���5=���2z�W�uI"DlM8�>-KP�dX~{�aZ.�ԯom��	H��|������<|.$l���X��p>U��F'���:a��,�=
RZ�Y��k����O<���ij0����#"F��I>m����[/��6w.�e�������Q�GfX�A.�j��x���W"Ů�N�'ܟ�Y*>���Џ����|B!uy��$��$����kzKc\��2$z�B���;P�N��q�5�g��,J�7ؚgc�$�Nb�O�iR����i�_!��-�4Ќ�Ի{����nRt�Zq}�/tm� 7hkiw�8���#P��t8n��W�8G��X7Y����zOT�>���pK.�?���m�}qP��<>3��K����zߘ�R̽ ɰF�4mw���<��?��W�;�w���|E����D��*b)����B��P$BX�#j��{ ��# n�zP�0����;�j u��\�YL��7u\�����&��MZy-RXXlC��"�ih �����������s)ι�v�/J=���u+�H����D���.GZ�/��ئ���� ����LͿcG*"���Du%��Pjz�*���]g����j��c�1�U��T�����F`Ua�]���nՅ�'z�ɤ��u�����������^�l8z��@�綻�yf�jUUeRE��M�Z๣��Qt>�I�$4�e��G1����� �8y���l���w>�.��d P(��/w��ۗQ5��1���~9��v��N$Iwn<	1�>��K�����4�s���z��GP��OXx�v�~��/�x�H�(@W�;�	<��W�j{qT��BNt�/�:}U���ߪ�NNc�Ug���P3�b �b{#��a,�~Aր�W$�?�2�ԓ�R�N ��(��rÇҫw�ш�ʝ'[i�K����ٴx�QN�X�?��j"�_�f����gAᣟ2���A�B��&Ta*������>G����x�����.;�TeUDo#��n�U�rӾ��Ь_�8�\7�+�2��W���k��<��-�?ZZ�y����q
�	^����F���Z�}�vȂ����0�χ��(qZK��5�S?*����dGs�R���K�}Hef���vT���d^�]]=s�\���.f���7�Kof������O����Ѡ�k���i�&���~�[l��р�!��'�a�wc�-���9��G�:y���H�a���W>!�>o;-k/au�Ce�Zw`d��6�AhoW1$JH���H�x��JY[�i?�����L���J��ue�1����hzV���e�)��ML׈"(}y!�NC�)��IGپ~�_�� �/�Q=�)�_��c~a>�%����i�Q�_�3 ���GX7������!4�J6t�6\Z�7�}̨�h_r1S�}Zݣ8��yM�zL��4��d�w��=?��ʁf���t�3x��,/��/���D$!-�I�{��N .����}�,�fS��*�@��	6�em^��H��̕�1�:g����
��NECJU�(���p��݁"7���Cޑ_�ЌAG��RH6j��x�-7q������d�}�@��Ś�
��*�A��[b޲�'��N쫇�R?QB.�`��)��Gcx8�o����Ț�i*Pn�a>�����*����"2K�y5��$�C`	����B�)�ZK�������w>K�<�����i�|չ�2�{IJ~S��U�ť�`���(1NV��
`h�ndbE`
-��\3&;�YM���c��w\�$}��'��1�Rհ�h�2	���ш����z�4�%Pϕ���l�!V&X=�H1ji���8 s�uشϖ��k;��\H�6����btu�̒��g��ώjA>�3�ا{�r���t˰�[+L3dېq��c=���l㹆�W� `Ȳ������g�^P�h��BA�U���T�]��-������0��f��57ƁEp�t���	_&��p����ʗ[|e��kM�k�Tw�K���Y�ҝhgϨy8�nj�p�t-?�%���#���@���k_�����Gĥy��7��+J����B�v�@��>ȭ�*X�l	�2�> ���Ζ�W♂���罎/���+�G���Rњ��L�)삢FFc��8)�S�E�Y;,�TQ�S�v�7<'��$�� ��g�$>���R�X����������pr�0�������z �Y�{��a���de�`l�n�0�CI�%'�{O�#�^�Y��!�N��]H�B�&lՆ�O�9��-X"�²�����2���o���^ҝipe|�`�G�#P��`�1k�m%d�H�����ࢤN�/IM�>��6,e��`}��ORG�d>{��!��0�	��"�$w��&kA���҈ޥ;L��]��l�D�*���� p[g�ǍI&` �\��?�}:X�n�M���>�I/}��~��}\���:��ɬj;rDI�55/NT�4�/J�25Vo
w�O���x#�a\{h������rھRL��q�F�_��+���=K��Z�!6W@h���S�r#YE&!z[-�f,�z�\�!�7�]
,��<�����F�a\u��x\�*��B7���v1���N(�E��jĥ0�I����'6�����R�J���P�3����_�{�L�B��ˢp�e����4�9mn�o$�>3��4�S�ԥ���1��� ��jһs�;�ߌ͒9�W��áC��|TfB�O�#�@TnF�sCV��y��������vř�E�-Hu�� ��]��)��|sɷb��;V�Lnn"z:n?r��]���VC_]4\���Τ�=��W����')i&}�����b��|儅��0D�k�Fy�������o�D� ��4�}b�TT�I�s���uj?r��:������W4:�`��I����H�'�b��_�x��޸k�7�7"���&��9�6�z,�����,u�}Pa4�s�A\�67kR�M�(u(�Y�G�à��t��eeg��g��)��������	��n�XP�����6\���R�r�����O�b~i����T���G �G����Z�#f�Z��%�|�c@H��������>�N8�Q�v��if3P$|H\�V����reb�
���(ϸg�N`c�X�਼ePZ�"��_��_�.�Fa�J��t2�uܺj�/}�<�,jfĹs���	�����MX���ȁ7�0G����L�{�<�y�]U��W�򻔞/�o�����oM��>�`�o�o��������A���~���Y��uK`�ܜs�e�Z��hk�'������uq�P��$=Ѯ5�A6c���~@�	�٩����]ŹjA�1/���^�/�g�����:���Gi؋@���cXy|�s��E׫�jQ��z���8&`�B��<,Z�����a)�I�t��J�??��%LBh�ws��~>��������_���D�88hV<̓�l9ۮ;y8$�x�V}A�]���?��jRt��lN���c3�݉�H����'�2��4��� ��[ ��ei�P�����N7u�r���F1��!n���qʋy/�,���'JGR8Gr�lA�5(@�b�*�+I���<�$vے/G;YK��70�P�Ͼj�a&2���S�?xxg#���@��_59�@@_���������������H�v���S�~�����nL#KY �Vf��w�rE��_���'��W|J�F-Krm�l�'����1P�`k_�Y��;�Tk2�T1K�l8Jɼ�d����q�R��x�YK$�58IF�˳xvv�T?î���0�@�F�z�y���F
��T�:	#]�$z5�;�=��x
Tf�y��|`;�����V�8�PK�Iaa��0y)-s&��6aֻl��]~�ܝ?<B���`�!����^{:���}͌v�	W���L�����LzޠL����W��H��]���"��IN,�}�����U���8QR(q wp�Y��'�*n�`?���FqдRr��$'�l��&������F�scf�u�%���Y>�J���x�Jf`��;��>>QU��UvGL�3��'��p�Io�p���GV$�`a�?�=`t�~��e+��4���0"��x�Yg<�����Z*k��'UsV��Q��CC,h��5�y0�;�XҝT��t�7�=|�}�0��w�7�����@�]��������m|������ 4?$�<�ٗ���t'����}%C@-NO6O> ^��Տ�*I���"�x�������Í&��|�M!�y���a���y_��/פ:9-N��:�̼^.%�����i��Q~�@�v�p�2Hb }�W"�Xg=P �=��p!�e8"�����H��U.�0;CiJ�3$`?Y��˻cM��[M��^��~zӇ;^`wAB}��p�21�{;��̧�Kl��7J�ǈ�a͖�N��B�o���ݸ�SRʺ/�*�|��� t��vUJ~��򵴏������V���m�}�-�]��ӿ�iyĕsf�e��k�8����j0C%�\@���Cꈮ��Y�l��5½5=0�3��b���Ws/����H�mzmH]�ɨ �$LF�����b}�f2�q�˱�+���2p)j�o�b��(�=E������8�@A��Pdq��۷S�����p7�����PgGFi�.��R�0��J�kW*�Ԡ{��mt�0�b��]b$�����L(�����tzA�ekv����HΨ�5TP(�	؊����'�b녔9Cne�Wp�w��=�*r��k���]���b��>��t5��R��z��j��&m5CD�lv��Ù���7o�L�kƩ9/���;�K�t�3=�"`�����K���b�����F�vx���[:k�!WO� �)�,F86mY���u�c'��~OgT�/��,iq{�ۢZ/��Rkz ̀����BQ�$,k����N~�4b{bc[Z�Pg��~(A�W�AI�(I���Q6L�`��J�R�pvEꝈKlT�_��c��:����&��k`�zƐe�������M����A#)y�罊Ì�Ն@�D����vC���鶳,#P)y��1μ�˰:�x�A� :����zqv���bf�EMc��TQ�cN�η��=S��Ec %�*Pr^��;E�����5
�s=�b�f������F�YqC9}�`��������?�%��Ϯ������z�k��-��O�oQ�4�t��*zһ.���t�ж�Q�$:�߻!N��e�G��$^�[�n�!�W��C.,?��	���)�h�Tr-f']5s|W�p	ԝV������;�PY�0'��Z��%��o�tR�u$N Ǹr����h\ʒ+ß&��v`��Lݯ �12�٢��[�m�!H��[��m9W�ψ;�����~+ض�^��,%;-1 Ӡ�EִЪ�B��2�=F�KS���ՙ���`%��p/��)ɏ-n3
�5|��O��LLLX��UϧG
O���e	��
��x�J���
�W�
�x0}�T8n#B�H�_c�d��LP��6�תF{I
v�"8sr� E�h����U����sX��r�Dm���}^��F�ڭ��ѝ1Ѝ��#��˘�:r����J`��Õ�ֹǢ3"���C�S.h]������1s�)����7y�����A~�ATUm5ݢ�'�>-���Hß� kʾ�F�(��������R����c�2�1�k֥k�<"g������6�|=^�HN�H��,)h��A�r�I�R>%!��p-u�����L�(��M_}�o}�͡�?�́��~\�� T��?f��}V�:���nk����
����K7ɦ^	�����������ѿ�	W�`]���Mo3���7�'Wm�3jQ:�Ю��њY�R�G8c�)V4@�31S+�ғr�z�n��.�5���f�u�c�����/�Ndrk	s{��;� �p/~j��#�%ϫL�۬�+Kg�cT�/`6v�����xl��̉��*Y�M�Qh�䠪0����=6r3�=�i�E������Vmp� +��B^8#{�ٮ�fZY�S��'8������k@�G¸ÌG�E�I���lӫ��ck�A����S|pId�"�b�w9) �$y�d��e@��W���^Kɯ#�p�Q}y��a_�{�g�vv5�"���񆢌��vY�������l�8�(K5��|d�&���1]>�M�؊����&����fyJ$��U�!��p�#��m�*2�~��(��r���P�e'$�դkP�uH�a2l�G{�4�G�9Ѵ�e�4��]
�6�*h"�����Q�I;h�\<�z ���TV`��;P�2�Έ;[��s4���"��N��cG���xU��a#��	�-�˺��Ҁፚ�?'�����c�n�A���pK��ig�����p�e:��)0;D��d�מ>BҖ�e���J@��YB��Kd��(�K�}@	+�KMk<ϩ� l���F�)�\0�e��=��oP���OA�O��q6㩈d�:.`Έ�/�)k)�� ����uD�vs��Tz�(e'L�?����XRm!��7�P��%�Pnr��x��p�����ѲG�3$�� ��7a�Pe�zv�e��rJZ@�@���>�'r��üT+Z)��mp%4�6�����	v��D���H�\2�u5��* k��>/P�I���/��_ݗ�*ƊM:�Ų�n�:I7)��V�Se���4��)�K]W�4�e&��aStH ����7�<������w�$}G��#4|QL)D�'q�S!����b¸���=�eΘ �� ����0�čW�[[Y����#t��%7��2\� ����N��9�*60�*�h6��A����I��2���+wh79�#MhOm����Y&������߾�t/6�����U<���j�e�����)�qJ�A2�3a�E�A��&~��7�;w�����iVg��8�VdT-zӦ��0heMڒ�	6�z���4��qm�{����-��[�ő�Ԯ���0{e���� �aZ~�+'�p��[����^�ZST'"+i�8I�p���q}i��n�gϔ�`��,ۢ8E���i�f!ԖtgԪ �#���Zn�!-]sӪB=+�̤U�6��i��(�Qw~|6�Y�?��l˿P��+��dR�=	Q4�%�kH܊��A&VLB/���_�s(^�6�!]�i����Љ��`����Sj��I_b�f�����-���:��b���$0�K�ר_�n��ˤpp����T�O�3nc%�)�b`�����\��o���������
���^����PL�W�^��T�!,r��U1��G�1�_fB��d�S@�`%".���fϋ�~X�4�Y؟��W\ǣG�4�i����v8�7�K��갓�My�O��	z�$�e�E��.�cꑗ�R�WxX��3��mgDJ�����ʴ�W�<CKŶ"xR�*g���/�ktB#	>''�c��Td�I7��Aإ3����	�'�ٺC�,ߑ��Ig����3UPE���?r����|����{[���l�ɯ���Vp^B+U��ej'/]��"%6ǥ�+��F�٧���gЯ��$�wy��^�~���#�?��F��z�)x��!h���'�C����^���b�p*w�(q�S��:�PA78#W��¤c����Ji'&Υk���h3�+���:P���/(�XM�Is.���R�y����<y�v7`��+����ղT �HdfD��!{���$LLb�m���V%T�%V��y�A~����?��i%aP#���\(D��VA��'��i�w�]�;��q�@�#)��w�e��k��Wn� d��\{�o�A2804a��yٜ͐�T��:����~Bs�$9g ���E�-�@΄�e�f]{�]�W�Pn�B�Z�@��Z+	����Q(�]���k����斊�S�y�Il�B��m �<�*,lKl	eb����cW`Gj�6x��q��?I�N2 ����G�&�!��O�o�<��r�6$�|$K�a����Z��{�0��-2a*��l��y�RIQ��%dI䣢Z	������(����kKv�B�*y��`�Zy�4|5;&'e��/�.�
�H7[�I�.�,� ��)���M����d(���7U�ݞ��DEZRW��$���Wֱ��+�ۂ���d�+�$^I���d��9M(�ӈ�B\�hm�w�3긒|Yۮ�7����#�[����ĸR�d����09�k��d�����E���{�>pݘ��i6�B�b����*���f.��1��NL�nL�cF>�A���U}Ir�sR�䗪/[�SR]p���ыp�;U%h/�<�{�͕�n)X����`HO ���2���+���V�2�@)V�c�P�]F������`jΨ/ˑ�f�AV�(>�g�H>C�+�d'�ͩ������oHD�UT�6 ���i���ϵG�03G1�3��FX��|hݲ^��@�������U��-����\�C�z�C�'6�߅�z'�@G�t(N���X��]�/DQѦ�M)������Я�#c���b�CR�o�忓q�ʖ]�vd�l<Y�������c�J/��s�l�G*N�ϣ>��W�N	�[�P�z�}R�cc�b�&�&�'y�,Ҳ�w_�hS�����&���Q��Vs�� F�ϿFSw��/EU���z���q0gxH�V.���z�H,!��?��1ۙ]�Xu���<��!/�����mw����&Z�}������ 3%���b-���>�<"Z�4��&6���mUJм.>�1تX�Q���R,`���|P���^Qx����/�	:*]G��E]�V�:1<���
J��M�8#Ex�`����F�CI`� ��{��6Z�G�r�C\����������ۣ�0��j��+)��$X��,$r�I�ǖ�@~A��Ně�-��2ѽr³j�D\�CΕ��ؗ ^���� ��d��Ď0�*��@�[��g�fA��8��x��O�Pw����?��|�{�Ue&a(4���R�8A��Aٻ,�n��"�
ieX�*�F|�sױ���ڇ}�x����j��2�)vP���C"�y/<����YD&��~"�����v��h?�'p���>U�wn� ���^�!
�S��T5n
Y)��A�⿉����]��)�tR����u����H��w�{]jp�7��hڇ}t��ӹ=�R�� K�\��!����M� &s�BƩ�B<[�������Y��׉R�0�x`3d��/�o�S�zA���Ge��[����S���*�Mb�Xs�>���٭�|~8��|?��AP>�Cv�i��bfI8��1e[��l?��J��n��+:;�@���4���fS��0{�s�%�)7�LT"6H�h��!���%wվ�O��^@�*��TU||�7bs��
1ޫҿ�z�U��yf���f�`6���}��vˎMľ�c������/�j��p��k�����~4hL�`�l��4�Zd���~�I��J����?�0Y���ב1�lܬ(wb����� �n����:�o*4�GX9���|�6��D�F�Xx S�VcG�b�n�$�9F�JsT��tSb�+�1"`_�@�Q�~�tT>T�E���L���чIv�H�G����%]�Z�<ޙ��D� H��QC�T/'I\W�5�Q��e��?DCQ�gM�/dSfo1��'b9nZ��(���*��.~i�z����al��	�A���
Yp��B�bT�D�����E�l����Y�/]� ���TtH����"Q�]�3wBQM�&Oi��\���]L[��;�8v����p�cĄ�l�s̎��9�"�o�����������i�+�����Da$Z�Q�ip5ͅ���N�����זPՍ�*m���%V����>(�����לT���jF�y�(��bS�Ps�s�^� {��k"�V�����B+�i��:.���|���Tߨ�0ѹ��"�����'rB�igt�|W?B�y=�g[�8����b��Ji�
��A&[��p�J��	g�5p��":����뀄��v��������f�B4N[���8�H(���|T�BلΝ9]���J����)�c�S�E�4n�}:�}�zr �Q�A��^�ӱa��F��Js�-�ƌ�%t�zMmS�?��U<�R�~K���`�����h�γ���S��&�9S�2�v�T�"�_/�y�3�:0�.cB*�x���9�׼6�� 4k����~�u)H&��AD��'�T�?Ϗ��"�a:��ɖm�֢v<m�-�1'�9{�^b;K��c�}]�����Y'+�Cvd�%l$�@z�T��X���'~���M	q��Q��A0�4��I#��>H��듼��8�R�S�-Z=�!:����*ߡ�:y(��*���آrtt]���B��I%rF��Ǌ���NW�n�"r'���Ov#=t2�\�K�> �蕞��'q!֌�x���(�8��oq� �N��FJ-��#)ۧ���>^"͚�k�"\ܺ_)U^E��ƖE�M�q�I�fؘ���T�|��#��k�½\[l]�:��ڎ�"Ɲ��>4S��l�vK�Ln9�j����2Yr����F�9�0D�]�;gP&{s�ۣ&����B�
�^���u�sY�Y#Kj�t�Ag��D��pB`,�:���K%�6��^��xP�\�Cw9·	Ѻ�"�qt�?�f�rf�����I\l A�G�ʡ�m	#-��;2��N�.���W�Gs�儁ܔY�~�I�č+Q��<�I^e��;D���I�������x��A皜c���T=$������I��_�J�CO$]^�&#� �DOyN�/\����H>T҇Ek�9�@�q,��C�uS���ӳ���:۪���j=�˒$Qi�eT�ߘΑ���8}�zFV�d��8�x��v�;�uKT�9��0&M&��Ļ-u!d%�8*˳HA�b�~��8&'��-3U/]��Z5�M���T�7���m�#!���q^��N��y�D����rD��F!?�K!���:Mi;O�#�
9V =��]����M ���LV��,�6&�,�n�^�bse*tCһ'�N9�`���\ ��m�*�&.5e�U�����Y
)�����P�3�f��7�2w�,��O�J�r�C`_��w�W9�n2G���6�����\��@N�񘸪0kTq�3��Y1�H,n�!fʔ!�����*2�]�# ��\��e�'�V�]M6��@!V��h�϶���O%h�QI)&�.��t�$��}H��:�{��ӈ�s��*�J��M�M�}�*r����L&�ȣB�l�S� ��V�zO%!��Y�p\�UBnG������P)��cK�o˽DZ[�b�t��!!���LY�9������ ���ǵ��pF�E�9-=���2x�`� 6QqR�8�9��Ǡ�1r;T�����R^bE,����~�N�L:X���v���M�;9�ϟ$���Ȑ���qi��?I�f����A��\?q1w8J�v��h��`�n~ga�+���
���p��l!u��q*�L�[@�h	I�쐒>�����g-0�?�#m/�N�K�~���x�Lw���X����ȧ109�;�v�@���ǩ���cT�@-c�,4\`��R�-ߎ������4ee�Ȑ���A�x�����3KuYdCkZ>�Uv%��$/�3��tQ���r|̥j�'c�
�[%-����
pv
�xg�{���>��?��kJ��#)jha�i0B��tɎ���HѪ�rL?ĄU���:3|�����p;�������<���^�>�s͵?�[
bݘh�:rqG��I>̕U=�z��^�`����<�?g�/�{w����fJ��M#�����9i����$��͝�N)):��ܺo)�~��[�Es����:�\��t�At�"͚��i��0�"��P`L��Ŗ��Q
�+�<�4ߏ�Q��4(yJ!���x�1�篘�������
�^w��!�Cô�yN>d�b�<l_��z^_^!.N1^����'Q�2����M@���3䃾�?�ڷ�Tw{�!�c���ҵ��TbD2�+�Re���b1��In�� 3��U[���v�Щ�����A��n�;�[�
�Ϥ[�@͙���x|�ܲ���E@q�a"�$5F"�";*�	�g���R��ZN����hF-��rQ6ZUzw[����}�j�����e�C�4L6��]��A�a,��$�e�%��.���t�_{#����2��~�SQu]�H�u�F-���g�8oc���?�����@��>T�A���A/�����8-'���|䮷�e�tw;O�
�y�E���|�W�+tD@\���p���F��[��U�xgK{���|�Pu����<�|jf��]���h&~&��T�rKv��_�����k�0oj.��0��䔜���y;�e�'qf,�c��ԃe���+��w�����B�n��kJu�pj}_7?��q�b��䨔_�x���#S\�G�҇��	�!�.����_޹˂W�Zw0���)�J�a�ȉ����	z��K�u/窶�L�fj���BdI��h,��{���gDW�.���ӗIAj�������1!��K)�>��^�P4��/����Dq��7�O�*8i�]�E�j`����@�Үl����̀�\֝3c����w�O�iD%{Qh�h��[00�y����@_\����$�����+���A�e���>���H���=��i�r!���m�_Z�)P3'�Y�_�bD���x��'f�g0�� ���+�!\A��1���R�����,��
"wK��?�+�:K��Ń*.��p���:�U�ՙ5��Z��V�.�������*��#��黹�؋?�l\:��^�(5�u>ꓤt�U��[��m0<���^��a�+n��_ϖ�>��,�H�[i
P-�Z���v�ef��C#}YN���7N�f��M���	��:��Ҧv��(�ك?�1�>!��l
�ҬG� ��b�+��΀��w��t9�O�lQڭZ�BH��u
�N����ۄ|ޤ�L!y�M6��qM@&T��&	�W��P�����'�d��5x\��O���������a:��]��g/u���,jx�SF>��r�?T���ʁ�h[�|5Ts���
y�ς:m�20jhI{&���G�i�γ��0�<%b`�U����`u�	:��Z~�λ�fjC�7�uQ;�HTZ�W���N!����~�ME�dX��K�=��񅇣�m�����*�������,n�o1�ZŇ�P��^����������A@{�;F��3��'�X
z��9;�2�ĝ��]<�zw�92�����@F�?te���r�"�(�p �o\�7��	\��e�{&4�qM�[,ٕ��'�
J�Ҋ��:���)��6�=7=��8���`���>VA���ʛI�P/�;x9/�qt�����ީ[���6a-�V�A�p�1�E9���3�m=X��`�����<Q}sZ��d���xm�� �5�q�e..����P6�7"�d���>��.�|��'��ۦ����!�y�2;��(�'W!�mE.������c�O�˺�wgƳ����Ve��Z~H�hh�~�[���.K�M�������z�x#79���*1�:.�#��'���8�1��s���`>����^�����t��j|`Aiqæ^'>�`�H�3�٬��w������.�pG=�%��~��e	ypG1�$}GyA�KLX4��@?��h�q]����kN~��iA���u6r�6ל���5�g����>�/��L�I4�@�,s�B�~�;�7��s[�4��10X��Ī�<z�����(���hR	���n;�9�ɋ��~�/aY*����TT��`��:�wHa��*t�- ù��ݪ� 	� e]������e%g���;�A-E˕��.L7�W�S�%��?�?��Cpt��|H��_l��I�z,��z� ���c��OP�o�s��\1&9��í�/o�����Wf�Fz�F����*��1�\�V3�)��H9���WǞ���@�;��	���9��<:��10�䲳ը�T��rKG#W�|��9e"�_�;7[g���� y~@Z�P�36�P��..���`q���	%ˬ4�׉����g(}
�$>i����݄�����^����G���d�b��:B�ý�P�]����PrX���#�N�V�IH�Qet6؄}G��a��;D����vc��T������d��~�xi�H��ص���]=i�L2;�<�K���+��UP�$^� Ϧ�
s�-ۧ��A����&�p�����H>�~��6�
s2㼨���"�{g�B���!t���@���_B��`A+�ݪ
Q�uƫ�ʎ�O����V��{'4��h�B-��-�߸שi\ӨK1pP��	tx��X�����M�'��1?��`yUm�U�m��JA��q��|�/鳼z�N�]�V��D�_!5�C�f
n��B�:[7,��=(���&��)�c�����e49�`������Y��˙��?���ȇ��~u&u��g`�$��>��ډ���������ס[��<00jOI.��J������?O{���A�D�o�	!Ef��i҉��gH��0E�
�RZgO9XZ�}5���o38,�y�E��.����"��>�V@(���f+���B����D��X���>;zT~��[�K�S�Ȟ�M�ZE_��ߦ���>�渜c֓��J���\�D���m?���Rؑ�=�)1�Qy11b��eu�Ӈ�~�2Qk���z��D�뙧�wLRTyg�����+}b�j��3'iD�z�Q�L�BW��#7��;��zr�t\�=o��w�)-s��˕�@�?:�|�Y�T��h��&.�5�#�;��O�4c�$E�� ͇���ǌ2Uuav�XRX�!ͼ=@#��J��f*ʉ[�a	��H֝d�����
d�Qc�{�K�+ٌ_ҌY-N�S�Ԥ>S#��t���)v�Ď��T��W~1)�	�QZ�h�+��g
8��[T^߼�C-��R�e��<�+����BotΛڱ�Ǔ��p�; ��IY��x"�@>���l�qo^Ř l}%&���������,��=b�18�ªu��=�l��q����ȥ������zpv�OD��v�,c��"�[M4�*]�eO��	���;0���"�@��ߧ�É}�� ���=�3H,.�ըq �~�v��͐P42��&�ZC؎l���A�44cdV��N4fን�b�HW�>�_��&�/�UF��n �8��4�+<�>���wW
�"���v�L��D�B<�2$�b��5�Q5̯)%ٝk�pƙ[��i�Qb=|�������V�|�NA�6���
w�� ���8��7I�l��w3���o�b����n��ҍ�ά�o�

Y�v�� )��p��$�P�RF�γ�W��q�	����I�#N�r�F�|SU��54C���EMH�?m�	Lږ��%�9�Pu�	�q/7�T�v�|R����^��Uչ�TΗʃ�00B!.��Y��T"E�z"Ƀ�yb�-��b5�w���~�>)x�b]� ̃%c��lc�j�B����<�-K���Z���!27}ow�s��@�6�J�����C�d2��L5�� ֥�&����y]M'f�[�ݘO�tq��Ŏ� 2�2O֠d,��[\Цu4�Ҩ+���)0��MًU��^{��	M"iu=i,�H:��w�M�u�`�O�-J����/Z�ӼXf�eK��+\_h:Is D�;�$��;�%?�İ�`��qN���w�Yᴑ�;?�,���mG:C��j�O��ʝ �1X��4mB�p!>���P��T� ��-��g�+Wk��]����/A��&M�?�z(���kh!:bLY�"�A�N#��D����B{aa�Cg����� ��E��DןW�]������u��LV��2m�n�]ן��Mρmp�uǦ͔-�P�=Q�A��tI������g��-Ƭ4!F�:]��Ys`�$�K���|l��A�@�H?F�����d��|W �-eh�a{m�y�{�vd�9�e�ѯ��+�<�$�_�B���٢��д�ѕsF����:����;s�%��]��9�檸��Na�̶L��i�*��Ҏ�?�����X2p�� ��� ���h�[�>�����hËf ��}�˓���M��k�2�j�g0�zJp{����Dl��婑�A���@��� o�e��
Z�[:��q��O��H-gf�d*��ha9��fÿ���B-<uK��x����g99��t��b�塽�7���zPn�X�EvH��<(�����d�.�#|�.��������L�_e��Ք�
�Zc/�Ͷ��
�bp�W����m����d7\�%�J����Z� NFQ
�+�������k�D�D�G�-��,b�æ+1��+�6�X!!�F��h����ҕ�� �LV/*ԀJ��'��	�U�Y������$�j����[�]E�t0�"�;�ў)W[�cI�����][ t��%�PvM"J�|�F ��J	�n��������bD�S�	�K�\��6G��u%h�6��8�T|��/w��:���h�fm��!󴛹J)��J��i�!߃^�g,E��G6�zei�bu�Y��}���ŕq�g5��KM��i�r��łN�؎aiRM��WQ���^�PҘm���DR���aZ���qoUZd�Sݠ�rL^����y:�["⥲�Ү�)��D�-�1�B��	��b��?{=A��̏d��6�	��;W��7�s/��ya]�'0$��e�ة��(ړ��Zֈ=T�����[�,#�j<>�=[������1x>�)+��m���a��ahP�눒�}q���G #�@^(�U(��z�u�'ɰH������i����r��[��F��3s3��vl�Y���I<�d�� ��u�F!-�	
W�-]��� �|]����	4T�ҙ�b�6��ٵ㥰B��cd��t�c��T�N��2?/�Vlɇ���Y�#��Q�iUL񔴷�Lh̖�ވh�3���EoN	���OEG�p����11%��bܪl��Xb�o��o��/K�����h����k`�Ӟ���?�}n���&y?�!`������ND�ލ�7Nܩ+Q[��x�v�)r�T(5R��n�%��~�8�6�C3��JA�Da��ŚN�A��O�^��w��`�!��^L��� �Y��hE�P�$z�/Բ0X��:%^����o���������c_���<k����/<�"����K<� �h��BJ���#;U?~���1*��Cp�5>r���>c�������t+J����B㲵�-,���.�i&*|�`N^��T�?����F\Lu��6�m^�����>�j.�jg�%ra�:�����cE� �0Q���Q�Y6	{M$x�M]*C���5��=�j�{�1'OzH\���v�X�'y�C��	]C���=�845}�:��(��s_h��1J��#h+,0��T)�/9%N*��[�aꜹ��Epm����b�[i;H��c���[�I�l��q��j�Ol@�.�M�P�B����|��"�?����3���+_�R掔�̨�`�J;0�8+�^o�̲8���(�_�����*;�dn��b%b�7@��[�ۧ&��-Y�d��(C�#��aJh��
ZE�L)mۄT��b���`ퟸ�9L�rl_|�)�����>�>���"X��w�2R\���B3JI���
��nr��5�̫o�T|ўZ������'��g+������]5Zd4qk����@Z���KC��Ɏ��hAr�>��0��u�<H�J6G�8�{QW
����& H��/?}Gp5ёp��T�Q�)0K|z*����h=�o�)�&V�d`���]\���?L;��k�8�h� Pȧs�y���o�iw��G�0 ��O?S�K�m�G����r/g��9���q�JZ3�\��0���3Ӳ�j�ީ�8�D������>���Z�$�,jj[y���IȣI|���b�̑���1��zF�d�[E�lr��7��@8�&>Vѱ.��6.����(">}��됒:�~���g��]�H�4�J�K���f=�@��O�6�����V���Їo�S {&���g$[�-�-ۨq������紉%j��vZb⊨M�����ޅ6�O���"��H��U������L�"	�ߩ�����s���'��i񛚥U�zӠ����U������@�hNʵI����ƅ�p�~�	I㰘`ޥ�.�B·;�Ǜ�x�g��������b��?n�d0�uD_
�ݥt�pd�O��1,]���y]����	C�L��������W���+dG0,��Ǽ�����)��ލj�3�����
��)�?8��{�<�d5~I9�8	�_��o�-B��v�\�0L+`���[�a��S���s�1��͉����륂��붗]�a��Mz2P%�E(��c1�U�V5��u#�ܠ#�ک���H�X����)`6�ޮ81ib)�y�ZcZd.nfRn����Fv�K��,�N���R 
/�����U����� @��高����Lф���^pL�G{�&�B��@Mz>�l2�O7з M�/P��D�膖�m�AZUd�C~@�,��mB�*��F���2�`Ę�G���ނ��1��B��R@Z[S"򉙐�|׽$�$˷~����zC��[vhF�eܯ�d%Ӕ7Nh���(S�|Љԫ�Zk��!�n�l�Yǜ����3�eќ��y�+�qHC��~�j�9\�w���S+��͔��RaX�ut��Xy���0��p]y^^,������^�_C(~���8�qk嵚�|}~E�!oZ(��/�W�@V.rM��C�u���J�:��¥康�}0�.��,��j&1t߳~_'/��y�N:&�P��;�N&�An#OO��֖򫬱� ��H�˻�z�`�F��/8;g2�]��Ƈ�Z��J��I���4_�ۼv�¼Ip%��L�oKU��=?��I[xN�'\N��P1���n�sM�]Q� t��x�ũ����ا��ݿ�!�L�1���!����ڶ�u܅\?�LW�ˁ8�����(�����]��u�y/&t H`��{᥍CZ�ۖ���NB�d��z�D�4���_�������X���E�{²o���'wd п+���:�p@	I�1��Z���ջ�i-�_� �:�2JHv���yȦ� Ⴚ~%�o��o�6d�0��x���M(w��G�����u=���97��>�(���_qNI���NMN���M 1�e�n��K5�9�s�׊q��~w�z�t�|8���-K�)ՂK3�5S�m�=o��=��}*\1�����`0F��UF�ۣ��E�>��Lk��A����2#�Ola�N�.A�m�M[-C��K����b��_}f�6��tB/�	�T���T6����{z�^-a4(.�f<i�#�]�N�-$@/���[ 
���:�K(�t
��}f�ioA3`$1�IK��b(8�(^U���.;W't�!X�k\-v�9��S����!��xK��/�'�hЎ5�jR�jh���6d�<uF������i�T��Q�-��h=����p�X�sd:�l�4$`1yu��N�}��ZU�l�����|d�S������7�Zn�6�vJ�߮�#/�Y�x�SD�cj	������	!��� �亽���
��bc0�,��oN4��{uAg�9����ԯ�w��e�ĳ,mL�]�q��m���I�e��Zq�=�32���M�@�z��Ej�K���Sjvl���΍�����ZJ�V�EVcXr%�({'����okܱU�����1?�{+&08�&P�3�y>PQ08{iU�-�0�N1���m���ථ�R�	Ō[�-�-9f��љ����r\����>�sv�hApFm�"s���,J_��}��e�qI�:��,�d�j!8�������"�|��8u�k�
<:h�~�6�M�8�24�{Ԏ^�6��Ehg�*p)�V���$	oY҄&���K?14!���������?P��3�BX�l�V��X�+��½�������HM��O����s�������P!��cP���뉳��æ8h��������`J�,�(}�q\6��_�raE�H2�t�s���?�V�x�0� �e<�y7�IZrzE�v�	��ގ��Ԑ�8)1rw�`�p�`RH�߿�9���M�^���/�`�����]M"?�%xi�&[�Ag�q|�u�$�L��3V�U0yf$I�A���@W�5Tó5�<�5��(�VR�%͒g
��>2vg+1��^�Z��]8��'�[	y��~J��NƦ �l��]}�ܭc�������d��~�C�>s��$g�@l����ԍ��}�N)R�T���[��0�uL4�|���gp��:nS'	Pk�R�y��>��֮�r���^ޜ�x���ts�|�]�k "E�ن��T���-=��ռ¢v؂V���� ~���t�y�a#��)¢�����]ߪ6����L�9��Ex�ު<�#�~z�#������r浞3\�i��{���4�N���!n���aƖ�yq��H,�./]��a�5�����Ȉ��Ҫc�4F�<�F����L6��7y�0�r6�W6���o
�����:P�2yg��&�!��#�!t�E�v(˺��Wh������R�|�2�~GT����'t��)B�[Z���n�����ut��
�F�����B,��0�1�v� �L�3�;�����hn���69+7���#�D�A��������&��BxK�ˌ�b��*�®��{��vr�� ����°�r�W�5R�OM��ڙ���t��#��15��ȥ�1Bj��t����,�Vbo�j�t�,F�v�(��&q��o�[��ׅY���:��c@��2E��M��e:Y���(����h1廱a�mf�*Q�d�k�g��+�I]�� I��;��3�/1+K�Q'�)7&Ƨ=1
|'�g)���/�a�1g����U���tk�,��z|_�'��EWݯ�*eɴL�B0َ���J��Nu�^���l#��d>K�"[>�W�J����jTĆ_�����|đ|`��z�&7�Y�Id�J�=0b}sz6�FW�6-ǚ3�4}����	s��2�6��Zia�p� A2�%���ՑV� ���Fv�e_ 2���s
��!d�5mK=.������~ԯ�`�m��x�7� ��};��j]��0�K̺i8I�U��஖|X�'	��~30�Q%�`�����fv���d�^�f�h��ωs1�<fJaa��W1�pU����v��A�i}��c�8��
P{�|@��q�����*ro���ET����>Εp��(�������l�jz �H1��P��>B�w/!��2��!�(ݴ����l��W�&L��Hx����r�� ��b<ؽ�bk����7C���!��j������T�ŀݟ��������آ�����^�x(�dd�T���Bv?������t,���+�}�z��z�\�3�"��m��h��a��MFٳVlO��Ɵ��9&EY�O�'�#!�c$(/���٪���l�E����~s�29>����-P���:ЉyM����"�&��=��ZZ��j�6.]�6�G0J���B��d�#K�*���m0f:<��@c�n� �E�z|���E����r$|#�e
I}�����*�t�,u���. ���$0T���LM����<*�#n|Uf���I��eV�ܫ5�˧6.�L�!~c���ԸB5_��sX�4�1(������B)�
��^36Jɧ��1��(6�Aǟ[��_�?ު���%RBT�G��2��1B��V����kM>�%�'B�����%�p�`���5�Eʹy��;����`����=�A󙹹
\4�t�Y�.Z�|<��n��&��A���ۗ苷�V�)�J��%�ح�N�`� Ij0�LZ�L�F���%`ؗ��  �uҒ��H,�n `jv�ؗ����̏��||@҅�q�r����;ieg���.E.7�t
6���	���Eq�P������&���VJ<5�g�|�{1��'?��,ĐQ)����|оW��ɞ��y8�᰽��X�IF�c׭8�u���F�`qv��ۉdl&G�
���J2������H���I:��\b�$ߠ��SS��Ҁ��b�PrM�(��";V�-4s<:��K�k4��i��<����@́��Ɨ\w�(�D��*Å��y�����;J0Q�Y_Y�91x��c�0����F8���D�#��XGvO���(���I��H��o$��S�6$H�x�1�1~�3�A,�y�����(!{~b^�8�NY�#������P�OG�������>r�!�})�T7RLPL;���b��Yw�M>��}�5��yj�=��S��<�ɩi�+OM~Y~���oT���N���k�|/,�F�c�N��'��v=���՞[s�EW���"s���d����b�����2JWS��m�r��;�n��<�A�BZ��bW���Y���>P��:�Skm��w��:Q|����.���o�"L�V���^�*	&��I�@2,%!6���5�~�z�wm//�(�-)�́��hy���47b��x� ��*�G��
���6�o�3�^��q�n�LF�:2@�ba��
qy5�p���t�g=�R�'V �k�y6���	Ʊ������!n/Q�V�;�2�s.�Ջ|�/%�H�X�9�`�MDW~(y�H.H�r^����������=�hA����.BH�*r�[����6��n���^2оh�s'�&��C
�n5�t5��Ll�v절[M��V^����v:�26
B̓�։��5,� ��$�[��F�Rk�22�ʮU"��iZ .��5���
�x��G��6��0��mWE��X����{��)Ӊ�C4o�Ɂ,c%߳�r�ͣXO�o�?/�>�hB~OL��L�=ŷr춨�`H�<��.�P�4��Ģ�x���$-��(2�Kw=����;"��:�G������o����.�7�s����S�Ş�@w�ͣ�׻-�w�ݜu2��R���e:��Q�� ��ٞ�!�t�'���gm�Kr|C�t���C��D��5B������t�w�0��b�I0��k�2��qќ6�ƌ�&#�>��r�����э��+q���<Qݑ�w�aqO�3I��ガ�b�潦�Y
1ɝoA �'J�o,���R%���@u��P�.�;�D`���
1�S�c(���O���?�lҷ(_�����X�M�'�n��*��ܵ�(z�z���-F!hͯ$(�m�0��ӏz�Cr:mBD�o�,�0g�����J,�&�}~���� ����? �#",ݙ�z��.l��-?�7���v�S����X�Z��)`�Ʒ�K��*�O��������VV�N��{�2 o.��Y�Â��V��5&pclyf�m,�Kf��`^��(��\X��`~��S�7X�R�,��h�~��s�Õ�;�W/hX����E�`�����"����A ���VD�POB��V<��%�9]QɶA����n�\�*�k~ż͂w
�3z�0��H06�|���0
Z3v�V!Q��
�GV��:w��啗��u�É<z���3{X��^��ku��<G3�WK+��"Xl�7c�z{��c�$�Cc�����[pwδ�V��7k%�ҝ�}�A�b� ;�.�M��J���"�p���p�ٞ�R%C�h�5Y��M}�`,�p�bjp��L�_P��Pa�IS�$�S<�H�W���B)�������?QE�ܿry`u�/[Utj	'��KG���>��T�I�k������4k Fp���þln-�=f�]���"�����a�F78ʆX�N|bH	��@s���ޢ�NJoT�J�q��xeo(��e�����|C(?JК9�Rk��6
/��8�>;N�]⏮�PK?ڿ����=�0�o�`����������2���%0-OA�嗵�YI�R&]F[b����i��}^�_��Ӹ�drp����t�;�ˀ]�5����~�Uמ��]*���YH���4�-�'�ۏ�qs=�6���Z5��'.�pz���T�%nGo�;�_zxa^O��[�EpaKq8C����Ll�+�k.r��RXl�SM�.�pO���M��D��Jܔ�al���i(����ʺ�I��A�$5��RI�fwR�Y�\0��g�����]g���7	�`��i>4<����=T�C��۳�YIh&�|�=�i����Jr���։(�!��.<����9bP'ga�!iT̋�ꆓ�<�F R8��q�`fxDe�;�ѓ)-aVtg�
Y��VE Ux�y�#�r�l��J�]҉��hX1�΃%�5��y1�I�ă��_����aG,��>˿�zp�Ð�O�o~8h�H���y&p-�ٴeG0g��k�ɵ[��z<_f%Ǻ����N��yQn�7�V�j�@�*�g&�t��2�`uv9"���E���	��m �+4'm��8m�xs��S��_�Rh9�Ҳ��]�M�)�D��v:C�p���]�Ξ��/2Ԧ�iׅ��	'1�J��NSbͪvK�J��$'s���N�n�i~�:�J�p�K:?;��
��e������4�����x�hw�/oƨu����#l�A��������G蛃c�ɑ��\5��i>�����NvE�^����c{p4ҫ�~�,��b�Z}�n��29zr�M�\6�x�v����:�'T�%��<��mZE���KS��j.;�jy'~�{�BRF���Q5\3`�@�h\�0>���������������:1��o�&�DR�	W�����9�w�&Puaz[p��lP�f�GSdVA��{r\%,t{��_�<�Gܰ��U���A�z~h�s{�# n-��̒LS�a�����o=��K�������w�[&�v�L�qﾴ�el�Bї�@OXrQ<}�u'��f�9V:Þ��R+����}�(���J'(��3�L�[1�|V���	��пU\h�Ϲ`*�E�3���] �������O�
.Vh^}7��/�}X�ۚ'"��~8+���H��)(��t��O�ض0����6�8B{��\�ؽ���۞7C/Z��T�o�����כ.J]^2��лraٲz��N�?����E�.w��-%����Q���j��
RϦ��|�����d=JvB��G�R�;�s:�썬/����C�Y*�GBE��@#��o}>�#�ӗL���E�^xnN����K[����x�a>8��y%j+*P���:�ퟻꉨ�B�������o��'1D��D풟�n��9\<��@��{~Cf<��aIc�l����wF��]�Ý��8r/Ц�w�HoFSK��c��ɢ4���ݾ���}M���K���f��0�7��9���mA=X���jL�|?�0ұpq����V�ҕM��D
l7��"�����A�[b-��� �kO��͡:�`0u��0��c7l�]26�V � !3`xe�۹5�e�[y�
��ne�ϋ��í�*�
�������l�G�L:1]���a\��lٚ �^p�)r�'D�Ć�0�"�b��Q���V}!��.�
�c��wP�q�0�O4ɵ
�i��>}�@5`�I�4Sk���O��?�����:��X�jt	˟��=�j��V�e"���	��d-^�E����چmai^cG{C��_��]"�}�JBD@2�ψ�����䵂,��z�?�@ ��+ڤ���k��A[$�$�����>�n1���]�������o�f�$bGq~�[?D�n�
f'�-3���'�9���c�p�Me�\�R�j��;;��ЖG�=���^�`�|gL*����7��jj9�e]*}q�����czY+C�S�P�牿�fg�j-�
���l��Ωv#�UQ��a�����H.��Jo \,��>�Q�I�m�ӿ��ԘĚ\�@_+�M��>���_O��?6�?��-ب���d�u
�R��X� G�������%C2L�k�KԙxV�ѼW��/�W·V&R�<�ZxS���}�C�,2�-�m'ᧁ��b �����!_X]�~���[CH?}G�Ѡ]�ټ)/FJ��Pt�2Q� �:�.�A'f�I+4�:��]� �5�H��σ�g�(V�/�6��+I<½��R�����8�����xs�a�l�`��B� �㮩ȴ�"�Y�Ϫ�ECM��p<	^���{X��E@�Ѹk�E�����M�181�A+tA����� �rOCk��d��zn��[��]�V��K�K!�8��Y5bH{!��HJY��C������,���~��l*˩&`B�U��a��w��T ѽ�(V�w�~]%{z�>Q������´�<�1P"&w?h���,���A�1<Y+������8��=��w2�cWQ
�W��J���"R���?�g�(���owE��d`�|ʨ�Q@�p�fKl8���z�m���C-L��ػ/��6�c5ӵӸz���J��)�J?��/��0i�E )����L���_e���X�"#g��$e.����T���ȌR=�N��7�1;$�Z�FPa���ia�ڐ���.̫��r#��c�Xret䬱�D+~���M��X�"��OPOx�/��vE܇�&EN@��m���
�-aVO5�w��0��0gPd�W���� T8�������}5�/em?.UK��λ����Ze�e�oT��(��;q�x��N��pl�"AxGV�#��B:�:�n��=]-7���s�{���N����\R�.R�х��*!p�8�߸ÿ����h��#��Z"�pn^��+cn�ņ}a���3Js� � ���|W5X8�P�wqA9]�Ӻ�bt5΁���*��x��V-p���ȋmO�B4U-�ڧ��f�b�^��78��#�z1d����Z���p�95Y�:5�U�"�@���	YM���JK�lGd�/��_��\� -�АO��nw��;P~Hڍ�x:�W*�_%�9�-�/����B�O�����ә}��+Ϋ
�B�\����������@XӘ�]⮁��T�����} ͩ��D t�^�5z�!͇�4�q.��耡�X��n=�K?P��Qb�o�쩪\1�Y��5Q�+\5tG�����E�)��l��Y �K>%��}u���J���J�y:w���(�̙}bR8o��T8���Q �lS٩Y"��$z�X�Zr|{���U�@�q�~�L��M'����%<�o�L�����k=0I�$8z�N�J"_�X�k�IB,/굒�d�XUq�at6?�)	�SJ�Ydk�Ox� j�� ���M�̜�����^��§I~�~ʦ��F��D��H��P�ɗđ��ה��2t���`�aI>��D���/�c�
��{sr��$�+��@�g���O���B�c�>ˀq�A|�%Y��:�-�F&.$�����`i^S�����=4�v���r8�X���ty�A�`�ʆ����'�p��5�	)��$�H�����rHw�����L�~�6!�$c� ,��[���$+���L|@�Wlu�m$Dk���6��u�g���Kh��p����\@�cQ����Mݓ��b�AaĠ-�y��O���ߜ�߲��a5��;Jz[~�+즊[�k����.`��nw�y�M�6�Ç�oY���a���1��ʜ��O"�ќ�%~.�W��d�H~7���DM)������>E$��4��L�b��9㐫u��v�F,b%��Hr^��Ȁ���_�0��O������җ�Q�h�C�Dic�������s�s����e�h���D�[J_|���4R��<��`�7\�����ю[�;w�4�r$R�������-ڱ3��ۖ $*�YI}7%z���3����9˺�u>�;)�KD:�a��j���(�%�E6k����~+��_�;�����ɜ��������kcQx���y��^�]]��b)����R:.ʄCvRH/Jq�..���gt���q2�3�Z��%���^HM%����<h�3���Ov3F�����nik�N�����f��/��zk�2"����I$�q��U���.������|�#���_�̻�KW��WKa�٤2���T-B>�_ipy��)�)ݲԘ��e�s̋�V�k�;�=���?�:��A7�E;Ͷ*�cJ�8m=��G�J9�j�֙��0<r��U�SR�(03g���*���[Aj�@�TAΘP�6͕4��`���I�㺀\�L��8T�%����xУ��\�]m�y{i��lR���$��1)�Ƞ��.5Q��}J������t
X�z-��K���S�cVY�
��|1�v��.���!2ގla����<�P��_?'D��o�􌻨��&_�޻M5-L�F{�k��fr�
k H0�c<�k��#��@�iХ1�l�Ǉ��qO� ����x#ZF���.��α��<m���er�.��U8�E��}�Anpl�ks��X�ˣ��H8�(x��E<�Y�ZJ��ǰ��XE�
�i��6�S�<l ��pL�KȣAi#s �UyU?�Jh�|@��B���m�7�F��]ݨ���i1B0G���"�������h��3K�AI$F��E1�a��NCˈ�����e�?
Rd|u7��Ȇ\���q�C�$�i۳���</���<^�>ˌ#2ڽ�w~�>�������i��uwv�}��l8'I:�ƒd�:�z��(���E&y".����ԡ�?[w@~�攪��>��X����FK�hYR���U++�����&b�@mt�_���UlǇw���kC6&Ԗ��Q$�R��I�믛g�0�9f���	J��Գ���9��%n�<H�#�k����ᷳ����M��2R(�J�&L���\>��?�yzxN�1��M��PV�u���$&���j�`7q��"p�YTl�=!d��?�J1�;l��%B	���c��G���eX+Om���3��xRG���"�#���>���a&V�2��"i8�'�6�j P.��X�Ո�|O��u�K�e/K�r��$E�@�2�Z��JJ����������V^�}�#��d���T�I��:����$q�>�	oڝ���`�ehW��&$��CD��z�җ)���q�a�,RF�����\ ��	܉�6��Z��:v�	���W����Ξ�(H�� z�{F�Swś�rjue�&Aľ�í+���2��|��M����X;/] ��+��0��}D:��3�Bs��
����G�l�lj�d]N���T�z
�K-ف6���k΋�<vVz.�b)��J�� �M�����a�,��S�Լ{tE��b�3i�����C���ξO��4�������B̼F��6%i~�O���Z���C[^�10�ʫ�/M�j�|쓚��>x������F4���z�bT���8��� ��l�e/]�F�u�FN@�3_BE`���J�OD<�g��}�u�q��� A�S�.���Y��6^e5 �0�B�������dTx�A��`�"�jj�c��ww�'L]:��Ė�t���t>�~d���N�ݱ�&\F�m��k�ʬ�;nG���l�r�N�K����k���@��WXzB[�8��?p�,lX�J^�u	�Xc�0�J��)N�Z�X�õE����z@���I0��e�Mʊ�g��;#�J��Yk�Л��uB��휬_��lѪH��ipp���g��T@���T�Vi+47����	�����0c��3�N>�b;���k��QRk+m��k�Spj��Q� �g|~��K?��	2�5IA��$D`{q�9�&�Z��18 XH�O(y$��(Bo���RX{��I�S팭�CH(O�>9y�x�HC�����)�cL�<�Ț'�T|��?�`#���[Q7��g���fgmc(�'�Z���EQ�o�y�������"�l-�Q2>IX����9�z��mm3M����Lz:}P���3�Q��u���l��G�7�q�5dT8��z�B�0P"����_�i�ʻϰ $=�Q�	C����*���6a�]?���	C��;�~f5]3�/����WGj�?��&�C̒��.����>u)~a~ �8)��V���%�������Ik}X�)�]�W����¥D�{c��s�X� ϐ��[2�*��<s�q�8�^D��2�ӻ�x3�]b��	�c���wA�E�]���(br'��k�e��������ƗiΨ����ۖݪ_�%|��xi���5�r*+d�`x����ގYV�yG[��֙�q���PK�ay[� "Ƞ�Nu{Ch�+�p�c�@�tNNR
��4|ݰX)漝&�2�@���|����o��ݵ�	���a`5lSW1ĩ���KW�A@�[z�Z#:/4�٤.���Հ�F�{�^N�W"YL����q�(G����T���Xٻ>�dD��M�qkz�*�2��/��ZtAS�����1,K��i�e�Y��Յ"�����؈w�Е�����\J.��]������l<����dg�p��)e�'�}��G#����ܣ-4761)f�_ֹg�� ����H:�ӣ����y����E���1۵,^�:�Sܢ4ht��R���5	�GR9*�ԥ�)�-�;�Yn����.���ྂ�U38�+Bkj���n}�6(slM[��Z�r���ѕ�yq��:�9�	ʨ������g"�>�_;b����Suĸ�<rYG��/�3�@�|�X+�m��#D���ȴ=ǭ�0O1�V���)��?��� �5Q���)�.K�=�j]��Bx-�!#V,�~��(b�4@�x�FAy폶��B��ӠO�Ho<�M$D�9Sx/�,t�u�_?(�('�~DM㛩��X���]ݖ&k�$�z�`�1�f��2��3��ɓ�(AS+��C�q�\��^�\��$�iщ��rV<�۟9f;3��*L���IB�M����ע�,�L��^V�GZ��|���߸~��w)<����;/�������\�p��a�i� ��9�x���,�����#�!3��
�UK�O��Gp��I6n�P
�BJ.�$}���tZ&�)��<e�6-�G���.�_e"��!�	YK��怂��w���x0ٓ+A�^Җ3�G����La�6��Ƭ�{�ƻ;(���?����_+�� ]�L;P�$���5��5�#���ݪH
�J�ۯ�r��Q�����`���Gw��Y�e>t�݂��B��hI��Ƚ�#^̤/.��	�ܐ�c��S�s�mY��]4A��o�M����Irx>���S�# ��|K�̪��Q5u� ��;;3B8�����������4%*��
�]$���wG�<�v`�0%
+�{��K��6�k��X��������S��$��XDQ8�= ��͎�Ew��ʳd�	��Ľ�j3(��::.���!4P���x�kSs��{��L�Kt�LZ�,�l�ZyQ*�$Y�X�?�픈�Ys|"�k�{�����O����>L���5�w�k���{w��O>Y��b�UD��*���a����c7�fif)ũ1�\���Q�Í����1'e���#4���#xD��ϳ:ә"�،d�3N� Ω�Zg&�M���(�zf��g1S�e��v��p��Ӣ/�`1f#�E��x��t3	�a��:
BEg3��ld�����Q@1��=u��I[�lblu����>F>#�|�k���[7]�O���/!䷳ZW�Ygy��\r�.��''���e�m�_�e��M��G׬~T��+��q¢��ʲ�������M�E	�݁[���<�� ���p�62��I����Mct���G��B9��0NID��C�n���&2l�\D82`dF��$J����W���aݞLy@�SЇ"u���D\��C���H?K��G`�a#�.���\���wkmQ�û���8.I��jL%(o�R_ ��`����G��1~V����դZ���KM�������*���H�9�?aOb@�f��B{s�a���������:�Zy ���O��΂�M��� !A�� �d? �d�c���ܻ�Y7��W֬���2�P	��v�Yh�U+��Y�	x&K�5EveO|/���碬��q�"���Jt��4IyWNhH��n�������GJ�D�FW͞ߦ�G0��~�c�������Zm�Ok���Ό؊L�&:�..���Z8w�a����^
�Ϟ�iF�%ED�	&�H'-/u?�x�� �'��P�ty���#�{l����h��m�p���Z�/v'��)��[;;�����)��2zd��<�I~��A���u�b���$��@�D�Jm��qVK9kB�M��t�Us�.I�g)c���<��D���:�[(nɧ��|54Qg�Q"��-���2
�+�Ǘ*c䍟�(����t%�	�*7�11 ���&�{�ZN�ǽx��ay��e�Ww
� ��#݀�e�*�9���8�d�l�C|WW��ټh��e3�d��t. {�8�!d�+s5�-K����U�{VNB�q|�I4��3�����Vе�`��� sy���
�\���H�]��h2��2�m���b,����K�{A]��Yb�;���4Z��
.Ѭs��U��%̓�`�$U��("�����:1,!'`'%r*K���\�%���^� �Ć����Ra�E�i_�L"�y>\�4[c���\�X���#�bX��.����{����R�� �5�`�ֲi��~�5��0��Ԑ\2^-��((]O��R�R�؞$��;/�O/2�s��'ՙ�^�ƾ����,y��'�Ƥ
�z_�6���<P��(Q=w�l��o�eF�_>��W�����"�(����y�i���< ����K� ��9:��@Q�R�%�w��[�2�)nc�f`J�Q��Csa�9�_Ӈgf]wfZR��
3&y︐dbu2��LGɠ��=0�Y�p'�e_�� ��w8�H�����k1�i�&W�c�ʼHRS��rtE8�B'�<���U��{j|���(��/�uZ���d��vJ��F��7����O��}����zLY��u�#5�{�Rg���
�=mm�o@3�4�c�$A�>>��׍�u�)��?v���E]�@�8wnj��/�<��`2��G������N+��ѹ�"�:�nZ���]�^#\���[�s_|}ݔ�֒����he�����P#d�,r,(�~I�|�(�"�'�v|1I�O�أ0c���x�yA��|͹���t�]��EL������c�koB�-���Qϊ ��%��w�Ƿ�L�m�O��iѳ-�f�-y�l��ZE�M�Y�Obʩ�g�"T�2�?��*6��dVq�RfE�c��-�y�IO�O4�L��]��Y�)��}����U���I�*_Z4�$g>�Z�^ʩ?EN���/͍�fdn��X��v�bxr����+���G�j�Y3AD�*�7|Ŋ'�N ��$��E'MD1��%v�_�$\��2��X���ːF2��ɷ��oo2�i��ך�����P�4���A��
9��S�>[�:n�o���@��{��.o-m	0[�VV=j�i]���IuO����[Et��1VT��G읪7���5R����Ag
d��l�>�xR1�B7�p���t��n�c��w��$��f��ە�\�x�����yj;�s���_�g.3�I (��"&{|����w�5fe;��qd [��U}��D�onW�bS7�ߋ��?P�����������%l��d��W�*N�	:��u ��i2(�U�hm�ݏ8���V�#Ҏ�>F>���9�hj�u.��Y��l��tS�7E�}���t�����_%�~uT��!�×c���q��&,�_��i�E�ݜ��=��BQAث��SY��N�w���Dm���a�M��[P���=آM�-��x��	iE����|��#է���:$�8����ʄ8 ,�#X�- �pwԮ%��̆��V΀�v�%ٳ﨓^73Sz o������Y��}���޽b�n�!��m�+�A�0k�p�*�aG����)����J_�3u�I9+��%��t����� �j�Gs쌚P=:i�3�l��-`!	'��*xo��Ͼ��5���[1�2�� ���6�9��@#^�Uڋa��x������*��@��WA8�����U���|Xu�h������	��/��*�H�e�zJ��Ց�"\�Irg��$�L&�ڼ�q>豉��ܕ�o�0*G��6u.졜.6kK�P	�g{Ɵx�S\�ǶZ�y�/�fu�8�]fl��+Ԙ��	J�I���gj(��SFz����b�x5���FP�,N~��=��A%��(@��/��dh՟�V��(�K:���Z��۫	�L>1s0�;`���+
�婍P���ʵ�b�8�c�����Z8<�KzU �z�������/��Rw��q�Z�X���D>�'}��sE���4Ww=�z������}��삪Rn��p(N#�~���1���Sn?9�v-������`���Ɋa�M�%���Gx6J-���Z����ʐ�޸���0�2-�X�S�C�!$WwZYEB6i�``�D����B��t%�.#��-�v� �تd��8(��oެ؀�{��Mہ"�d��tw)7�ٗ��@S&�b�\��m���ӽ:`3��>+䯷. ���"�����ZZ���N��
�����hSj.^�
� ���/y]��jR$�x���ls1V&oj��3�`B7����Xi����/�g������`�x�+��7B43W��Z��e�L�o%�gټr�Wp�.���Ou���I���e���T����n�aI �����:) ���HЊ����^q�٘�mQ@�!FڕX�r���w�5f,3E��s<���u�zA[� �����{ ��p筹�T���󦖔hq�zX*�Q��I\�W׽m����Pf�� -%�BҢ�ݨV����NI˨=�x�Ӎ�h-}����	�B`a��� j�|[�3A4{�N=瘤���h�"��;��l��s�5�b���	 4�pf�L�c�=�s���r�>r�7�M���wۓ�]��W�dv@�C��GZ?��[&�*f1�p�6=��ްqZ
�mi����y�~�ĝNA���J@:��I����/�BŐ^�,�0�rH�<5���[�]!c��d��g�G������7?쫋���L�x��C.e��QC_��T2�{&���{�;���F������柽x�?�S�������e���)������Hi�{����2u�H���5Z��$G1����-�����6cR�(8%3ҋ&��0�4�׈�i���A*�YA
?^0�Hp���H���
�ėɅb���ś�goW��[�
��_&�
F������ҕm�o�z$��V���;	Dd�sr�L�"��f&p��ٲ�١Ć�4�uȍ5I�cV)�_qOHS6����Wk�j�Ӊ��)���4��^>��ȭ Q�(�Q	��q��g�Y�#�j������͑����9D�l^��3�yO���EV�5~�zHA���l *�(��|I8�|=�V�m�B�}Iлyt��3d�����w��S��6e��הҹ�(ϕ��}"�
���o��N���w������1z:��m	��|�&e��<�.DT	h��w��B���?7Ű�mՋ��a�s�)7�ۙn;��M�	��d�Ӧ&��,5��ǯ5_���<���ȫ �/�1�3�n{��S+�P `�����w��`�=�n�cMI&^l����%W��Ϯ$K(��a����f 7�"2w��pځ��d��|-��ŀ,�_�81H�j���{>�o���+G�A����^���l��I��0��P��A9X�s)L��(@� lO)?�R�z�4и��:�f�����E.z��hV�AA��B'L=��d��z�K9'e�+��KK�&O���V����U��>�; �`�`c�Qe�tp��D���$3�^Z9��Q^z1U�#p#=�p6��}��)�t,�ƺ�Aeɇ
���#s:zQ�S�->������r� P2�ݮZ��3�N�a<���R�b=
V0�\pwo���
Iyy��|�(�a�TZv^ٴ�(��@իU4�T����G�qb{X�ؽ�@��v����ªԓaS�?PI}W �O�8��i�46�٣�M�t���bQ&�� t���7���˞�u�O��~��ql*S���55���߿@��7�� �*h������S�%����μ�F=�(�H�;T�B�A6s<�9���R%��[��o�P����p�"i)�r�A��
��`��x���́j���ˤ�bAcUן�\̒�9�5��;4x�Xu7n9�����G�Z����γ��X�9��n�c�gx1���Y��$�X������2Q�̈j�d�O���v⊧�����n��wѩ� �G� �����C�E��V��u!��D{���1g�0C��
�i�-,�e8�'蔂��,��Z���A���z7��3���l]�,�u]�5B/�J��s���|;�O,X�n�M�O+T����KQ����VT�������Դg�4pp�K�����b�V��%�S���hUu �p�����E*"kӲÏR>�����l��bN�Ĥ�Y>�����@>���uE��}.��������������_s�L2���[Ț��Yvl'e��oS�4���۝��1͌^1�ӐP��Y�k���u׉����#����zb�叩Ϛ��q����w|�r�QS�mRsB�`�ʛS�L�O5�4 _�Y,Ƣ&�Я�2��/ڷw�g�
����ߓ蕊:��I�W��+,�{b5s�_�.�7���
Q,�F5�E|ụNA�+g�m��~.E�m���s3��X��n����Ѭ�۾�ZO7��Т�bX$��X���Έ!�>J����\�-Ҷ8�,fx�+�z�5�q4��:�o��g4:~S��������J�n�r�#^�f�O�Τ=�9\0�1�	�"����>T5����.�$��07�Ho'k�L�����E8��3Ԫ��C����w�U'ݡF�/����(��J�ޙ�B�|e��Gǝ�MH�����y4��N, o��^D�f�ݐ��V�)$����c�fP�\�A�m�;�v�c;
*��H҉}����<��L��r�*�yz�?j�+^F�ki�)�ݩζ����-LNxG�Q)�+��Qo�!��%��᭲�Sr����al7_�Ī�K�0<�w�tʱP~�m1vUg�a� 6ۀ̦1E�?��[���=I[k�C�'.�<p��h����J����e�h[�����)J2.��2�5:�TS�ݟ�y6�d���(����n�F�<pD+Uck���ۺ۠�����ҴS�_�~϶"e�U��i��jO�+����@e%���>4���G��s�:~��:E!���ٕ	�b8T2���e�*�G��:�i�������|y���!ϥ�M:��!�1��Юie��D�c��ޱ���-l�K�T�s�:�١��l������is�=ol�3��v�������w�����h�	8?ψ3{���N�}���f $�b�Wu�t�GUmej7tC�r?U���>��|&*������E�v"����:r4�:/܅ͧ߮Et�3]�jw��#׼_ʴy𮋆iqs�C���K����M* �����(�����+}���jp�Z��q �4a���%/��#M�s�Е
07��KC�(�~�`�SX7M�9Ͳu����h����N�C��Sw�I'��Ű���;i�P)3)֌��WOCV~� ��59��4,�͟��V�6�Uy�[Gy��.��!�K�m\.M�kR��C�5��#L�ҧ�0�o�2{����\�mɧ>�Kv3��Q�T�^�o�Ժ�!�_���Ҿ�a	�+��D&Ǖ"��_�w�*)�k߃'��{����e�J!M����fH��b6O09v�$a��)�mX%�W�v��� �	gP����R[���9p�4��Wߩ��V��Ѵ")��ڡ�Bf�a���I��\��F�CBn�QBYyaD?hȄO���Q�hH���G$3�H�yJ[�6�E�P�^�$���!ӱ�� ��2����@G�Q�S�3E(�?H;	��v��·�*�(�M
�R�c�O�����������z��+w-��$#�� ��`�忆��]�,��%���)a�z3R�AY�ݪ�zqvlpR��UŏN�J��ZI��}攨��o�X���5���թf���Zf���DӀ��X>��������r��q\���S3P���6{���gJ.Yq8��f:�1��Y���WY�/g�ŎӤ�;�Jw�@*n�r�G���������4�H�E���p�~ox�7l�:����]�1�
ȝ��6�!���O�,q)��[l���ڮ� `��rAoF0��q�*�#vx�q-�ַl��ī�M�0�g����绛�G#���1̑�1X)�)=�XUn�5s��h�#R*�b���mH&DNvKBv{������&��N��D���e\��'0+�\ M^�㵭T�C?�q9���M�W��}&>P�B���i�"�Gn)#��1� �c�A��β������lC
f�4Xu�E+�`�	H�����(�� O�悥.=0��d?B�;�o�e�լ'��XU�-�9��J7��h�����YT��5������@g�&�����W�,m��)����w���A	s*d0�H�;Z�`l��t`��>�F�~tTɠe�~��rXL~����P7K���nǳ�\�q� ,�ʩ�7���� �ަ��J��&=0ФÂ�j�q,��Mፌ�w���UG%��a������ 9�с��U8cbi��z�|uM�J~O��qw��A[/���J��i�7�VB�z\t�i98�^:�ṵ́L�E�X:�ŷ�h���=�U$�A����r�uiK�G�,ꊚs麗%%�
�&��a��v�2%�N�J����SݴT Mz�E��c ���*�Քi�p��;k^#�U�0hB�c�$>�����L!	��7�+���QM�<�㘌�SC�AL��FO��8��D�='�p�ΕJ� ^u�xf����|�Y�o��@@f���l�I�LWH�8�)<�FjZAd�;��xJ\ozz^�Ŗ�J���� ��+�9v}���J_d��7��z�lpNo�>z$3�S�4��sS�l?t�^��d�$=����2�dv�#!�-h�$X!�.�[�������Z�X�+[�����N�Ҩ�Jwaa�ܒR�(Q�#���x�Ld���/��fC�t^\�B$	{����H��r�nS�c�f������L�T5�i��<�W��>�3��1(]���J���:qF��B<��6j~
��-��{��TW�"�L+�/έ����1��q{ޅ�\�[���m:H�K^�E
rV��3�������G��i�eq�	<�M�i�h��(����祮\��NYPT㇟�}_�U�y����e;��]�Њ=�{v������q2~�J�S#puf]����\ӉO�+�vL��c�;2��;�i�l��n�vܵ�����)0��Ih�#��ϛ��
�ݶ��J�g�"�϶��rc!��-}&c��}\�9�\iߊGk�7UV)MO�\n:�%潫1�h����*Z���;Dg)	],�B3�-�g��M��M���(ɴl���J��Q�'���Ϊ���^��g8M'���&���"��|��i�!3��ڈ�E��h���t�Iŭx#��:��:��4��5ڟ����� �n>O�@�9��.��^nV���9Z�Zxi�<��ÿOΘx\AMט�C��.��x^OV1�j�������2� [�q���'9�rS���/T���*w�ҙ��e�nA`%�Z.���� �)_�<�������2����0�g,�8j#�1|��__Y]��9�pvζ#Ȕ1۸�jcR��w3��s�E�J�~A��}3.BdW���)�]�m�SVF�(���O� ����"��R����6 3��"��tev�H"�D���-5ӧ�˞U!Q��L�� 1���N���bS�<ξ�����cˁ�]�9��.�M��� ��n�jQ�uR�70J�q���jfV�^=bM�!;%D��!Y��+4���bH0��u���ǰ1��*���L�;�ޭ�����bX�8���rAM�D�@�Oql�Y�D�d!������Y`J��8<+�' ]�~��SP%]s�9�'1�
	>�*�b7�f3Aͪ��`]�*�\��g��\~�V��"��*���'��|�}�n�A����mO�������#���������2���`��ɋ6�{�߾�i#(�:D��+� U��')s�T��9�zla��M�N�ha�"�:��#Ӳ�1����m�P��N��/n^InI:E��v�7�)AC��0�9�N�t���� 85^䣨�<k@ֆ7�㮘XXa^�$��^�6�0Z�Qb_�-��co�L��<���`�%��	���(V+h�L&XYZ }p���q�/~M��˝�0��b�)AA��S��0X��K=~P�%��7��+�����kNo�dEQ\�NIqX|��k��z�B�$Z9an�?5����q��FW�
�(Y�����?'��-oz��C(�6�d����X���5Y��/�LF�b�/Y���s��G#4M?��KP5�m?x�?#g0�=��ݩ�Eu��L�d�GHl0��y���\!�2���:¾�1j�GSU��v��|�
������{8aY�ƚ�)��ィ�,���qdHz3���:�o�jm�f�� �����q��N�A��z�ܼ���ǁ s ���*��n��쿡=,O�A�
��HG�FP�8��s�?®i�7]$T�f�l��_�sp�u�@_�'����i��]�*��*O*g�
.-c�z޽�HSk�7�������ݖv䊷XbeS�������%��Ӂ�Hv��L�+�_�s��K��.ɛ^S�ـ�n�:��2�%Z�Mݪ������Fz�B�������ʝi�cн�[���#;�1��eeڪ�[Ϙ��4��j��('�])h�F���.��xa5����ޛ��A��	��)(�_��"�Է:s��2�ʨ	x�F4���2�A�yL��6ܗ��=�l�+�[Ջ�N�:��ui%�@������J�3Srw��}�u�����h�h.!*��K�����Y�f�c�$>��'{O�æ}4�_�t&�t�6Ek�g[q
-��,�ObT��h	�������y��-z�,����}��N>o�p5��G���O�ޚ��Z��LY�8���'�+����K��嬒}3K��S��zA��u������ ���oq�����Q�7���S"��F��p�X��X�`�L�bi�]BYd<�A�0K`�˪8lDUY��^�7c�AP���4"�����Ɲ$�z
�%�����b?�)�[�M���c�=��r���"�1��i+�
�����)�M��;��%���X-�r�8&DB�i
����n��'Z--�ξ�E�t���Bh��(��D����rv� �]*�]��K��YE���˗�J��9�凱,��׋`�����褼�8��h��$|��)M��)T�b�[��
��ń��R!����+�ˤ�@���!�#�| g�J���4Ʌ������.P����XY���Ī����̴X�|z��?u�?�6��K�D��Pm4<Jĳ|�w78b�R�������7�j�,F�N+C�=�蕭@D�ji
H� �gH���7��Z��{���x� ܶv���[�C���0h�ɍ��@88�����s̩�(�o�xS����Ro8Z�����ܪa}~�
3�F��|%� ��4߭ˑ�Z�s���n�dz^�r�����N������v��/�+�Z��lg|�A�s�N�R���� ��{�y[�/���`=�Pᏼ�7D�zQL,X��g�U�<>$!>sne� 웂 e��x�U�=L�H�������41Zn�,"��&��{�v\$��ͣ��a�f �9?�F�������WJ%n4�폽�)8��3�e+!����xc纂p���ON��=l�.��j}}�bz�9w`�7r��dt�{�Mi����iU���фH��(�~�^yJ>�.e��Z^�Տ�B�	��׮�bFW�]+y!�9X��dT�\ފ�#�H��S��1�aܾ"�#J���.��^h��f�K*�*�~Qʾ-����O��zR��dhwjQ���SC�q^�A?�0��!��u�P�W%kd�T�=�Ԓ��4�TJ�.JJ���4-D\�؛F���=jOR�Â�B�{qoW��-���lĀީӍrm?�Rb��Jl[�ni����]�4��{��]}��!P�E۾:@�z������(
qN�&n~v�##?�J
I4'R�N`˱砪��aM��g8�}7][ZXKǝ�K>��#3"o��xgRVJeyG;(P�U;�cϳ��$��CL8�V�P�IY*���V�!aX�epURC�z���"��"";��F`(��ώ�{���mr��ĻG�*,��ђ�]݇�z[����n��&������ 1���������L��߂��{ף��S4&��f1�
���p%�n"�A��{i��ɘݹT��R�q��8}(��鞆>c_8���`B����0�ԋ���1�+#�[̘÷-&�Ⱦ��9�ì0�:���#�t�`*��hbͼv�R���h)<�P��jf�*�I'�D!�~�N����d.��b#y�w� ���|m���d��(��%k��ٲ�� �qM�剈��_�[ 4��	�",h��B��!P�f�p��.,��19 J��џ����/8�a��q+�Hi�O��D+\���֌.��Q*�σ�im�P�)�*�}H�P�sDafQ�.�>����m�?9�-8�+Z�w�c���NXL����Y2��,IY����Lo�`H6�I��q� Y��/�H��)q����y��h��t�(�|��b�Þ��~?A��	M���:)tfs�;%�"�����JJi��z��-p��ch'ч2�ݷ�w?�P�h�<�	g�h�/�o������'���8.Pp<v㴠|�uNlћk�~���Mk�;'��I�+!��l8=�.3����4T��}�\^�_G�x�&�:�&%`����(z�7�ԩ�|Ka�	�OcmO�����D5U�,|?�R��4Mtկ��1�r%��Nfa2I����A�)4s|x��o��4h���9�l8U�f�N����6��=]�44�ά 2q��M�!������<��NXɺ˜������ne��Eb���Y攮E�z��%Ѵ�pÏUGc1c9,����?�ۖ�wu����@�ö{��Z��g�Kn��e�G��]����9� ����uHPG :f�q�P;@��~�{�l)ːٵ\����)VR�Y�����O!��P�֒]������U}��UE���88����6��)MĿw�-T�B�<)�(��}�a��(k@&zk;�1���I)��K_�i���ˉW����G��(>v����^�b�'��z�!Mb�j��i�p�5j���_]��)�
?��32�yF����ʫ 1G.BR�u.B�)-Z(�:aK?LJQ+j-��j��)�����N����ۖ_�9.~C��������g����[����5l��o���w<���>	͑˅o�l�����ϼ�c(D��j��%;	�Z�~+B�tj����h�q�o����-��$�5����"��'�{&�T�ϛ�>�
��d��YA��"�|�����4i)��S�a�;ʽ�zٞ)ի�c���%R�S�� �?�4�NS�؛F�,6�P��6y���Ϛ�D��MND���Ӽ�y9S;Zԍ����ͩ�kِNo\�g,o�   "=��c��z�Z,���z�K��^J&21��@Dq���N;�p���~A`��E�
�J����SF �.���c��+$� �(����� ����-}x�̺���.@p�Q`}�F���>�(�(��t��8Y�zN�@H�k	+`��rE��~�w
�44Un^��ч@�x9:pqu}�VV����81 ��_Қ��x�Vx��G��T��&�W"�8<l�=ߡ��@6
��ueq����)m³�ฦN�����3��V%X��6Ŧ9��i� 0�D�)>�M��M�Ҏ�4�P6�^��}"�l��5���Ŷ��3p1n�,p��p#�L���0����5�G�e)\/b��w�fx�ؕ,ol�@�����/��џ�[��"Q<�������:���H�w�	��h&+ny����$�lg��ڱ�S"E�2���q@"Y7P�
k�) n�{DU�|��#��3}�l20��.j����l򊿊�0��ؤu�/�[`J�T�}�| r�7�wAv�ʸ�U[��o��,�%-��Ü李���^Kژ9��7�A7�#�ތ���X�w� X��S0L ���T��5��7��"�0��K��u7-�P�tL�u�$����eʞW�
r�o�Ǹ��t�w�|�xѤh�˓��͋����BN��ڙK/�"���l�1��4*�D�T2-�#Q��"9�d�q�\P��!$(g6#��]�ۅg	Hl�$d�:��3��`Js�V?/2�\W:DD����5���._�mx��b�	��;���~��WI�S��A��Yn̶!O&�#ܢ�!�[4�5�,8�=^��e���^�'Ry���D�|~Ĕ��$J�k!v�ԉ��9��%�3�g�s���Ľ���WM���HfED$�ɐ���L6����ӒX3��#��X�]Zy������`�pLZ�F�� ��}���ڹ]M�S���9J�WA@$ ʅ�E��A�l�1��Z���@޵FK�R
vÊ����?�a@��WR) ���?m��v}��̩(�kfcw�`�OJT?V脵��N�Ǩ�wr%��9R.���j�_K�*ܣ��x��-�=X����:��/�sC�p�5��\�+��ri��HJ��o�OU�d�A�����)����	��g�;_v	��<��ƣ�n�ex�ʀ�!jW?#�:L���'{iˋ�M~�*ᰘ���ḻS��hG�䛯	V�����$户���纋�V%���o���8�0�)Ok^�;����Χ�2��X��v�vjB�`��kp+���d��Ѷ��Z���b+-�=\f�q�rDp� Q+zRn�;L;?�N��a�Sh*�nĐ�%�Qx�<Й9�S������u�� Ξ�t�Q��#�-c�������[�̂�bSȳz]�ZL�h�=�FvMF(cGy%��B��^j�'�d�5������r��|�%��"����D}øLF�e�?��wưΚ�7GY��p�1�`~�>+a�%��W�V�<�Y���
b�'t2"�2sD��f��'J�G�ӫ}N\�[�꿭�U�d�&ˤ�$%+u���&�c�t������Pxev+�L4��%.~�^۩𧻓EF������t���qF:�E"fmtk�/_T$�J}�ig�i�P�<�HYU�������wv�Ձ��^����k�*��[1ṛ���ɡ?���YEޢ&���������9.j�*x��8XЛ�σ�\���3p$�;4�o�À\E~&�c�*ݿk����#�4e�Q�%ۢUA�g�!��:�e�K$��P�Kz��^d�%� �#��F4��q�D�� ���"��C:�� :$�>�d{�vC�.������	w�M��V�j�.�ٜM�"��&�$�i$z��'��/�����p�եnTF���f�j�|4���v"�	�iL��qz�b�d���z�(�X���3R��:C�S�TR�TI���w�"AH�g�����n��<���$�T��AC��r�a�������ۜ�������
����ܱ9>7�����"����3�o^��ȪU�u�?M�X.!����0H��3��,~�����������S|���?O(�QQ�a�r(��/�������|�d����p#⚶]�B��m-Y��C�Q�5�S��j��G�6�"�4~+c�q�CX�����oed�a���KS[Yro�k�
�ەB˅LƜkQ��_��5\H��l?
k�I|�>g4i���c�!O�%�����{�`�F]Uk�ݜ�Hǯ��a��h�r~���,��#C���5ln����A[[h2�C�m��5���O���x��N7���6`i�}�Ǎ��[lvӹl��V��ث������ο`����>d`sõ�>�A��z
B�h�q�8c��F��Ff���"w0�L���i�\�t�������d�+�sԤ���O0{vje��^q��[�gĸ���ѧ�L�7l�!�,�5+>�v���[������K�}���_�P9C�0�&:�A�#Y�$�ޕ�(t���5 ��t]�V�Hw����x��][�F���(��ހr�=�׵��`�)j�1�\p���J���U�y�8�*�r�O!�t6����v�0�8Z*��s|H����A�ꞗ���I���_H0�eh����X'��L�,��_�T�n����;G���P-+`�2�t2e3Oj�3���O�G$:C�K�ŤM[��07���^�=��:�cՏD�* ��e�2Ū�)]æ��刅���d�!m��W��D�"��X��0H�d��7�9�T �ۄ!k����>��щA��Z�+}� �u�����F��-�?}���Y�U�2��mª�ȓt��6e��;0.� \�D�0j��x��0������*�T���l��v�	�&��BI�$�a��?�h7:A�ᢻ~<�#��%��i�G���/s{\��Z,H^� �(�P�4�	Y�H2���xFSi���[P�R����ҝX~#�o����m7�PO���l�.��֠�b�w�ҋ��s/i�F?$䪦/�L��v[�ORX�� M��N���r�J5��Y���_t�3��[��$(
ً��WŖI�L?Zj�D��)�����g|�y7m�@�DA��x]S����/ݘw��_7���bt?ꖪ;��Lr����`���h��[�4fpX��/�ŜR+$w� ����K,�?�96V�v�`gb��3�>j|ۉ�mnp[t�		,�2ex����?{Т�3���s��`�%e��l0PGk�@��4ϐW��3]$� Y��i�s�$�|�^$��Kv��7b���ݐ�7NŐM���S��
Xk� �K�R:��$xz�2>�a�m�DX	z�"a�����ξ����
��bD�h��g�[��u¦��[��n�֟Na�����5�X��y�(�e�� ��7P�Z�txl#��y  :�H�����	�^H�]"���2�lY4�]'�+�xό�t��y���i#�J���q)H�F�K�%{�uɻ}vn����M�d!A�;��oB�l��aE�k6�?��ɑ��� �@��;vC��q7O�nHCWf�I��[Al:�}H�*5��"�ؗ��������� ���r{"��oCQۆ� 7t ���ȶ3��:Gޅ�a���x)��7�һ�q�Qrw�I>�"[�W)��3��MS�D��Kl&���֦z�����t�U3Q��N��\2�����5OO ps�vBg��
�aS{{so=��XX2ذ�[��}#7D)���u1Ȕ��O�N��
�<ׂ;����6�m�=�8��7���꜂�׵�ȏXg��5��`�h�F! �Wei�g=[i }�2>�r��wqW P��]Z���xL.�H����BGY�`-;�J4�Ǥ�ViZG>����7᪂�>	���!�9o"��$��
L�tuVr8Jg�<�^�aar�]94�ZNV�Zћ���;x�݂(��25r�a#n�p3H�\m�K��p�m�ľ��%|�����s}��LyB��;��,"P!���F/���5�1`c��;��7&@�����k��h�ӵ$�?��]�zn�8�?w}+��T'-5w�TW:O/1�{�����a�k(�TI���4����ʖS����)u����9����u�Snj兝v��2����%��v���25�Ɗ�*�HjWE2�_6$�C?裿�ڒ��/G:�{9��|1{|�g�3�]�f��溱i����R8��(쵘"�M���T�h�7C�I}%��PD�j	����t�l�"��W<�pn�p۹�/]�����[��A���6�_��ٜ�t_�Gi�k��=La����0ټ#de���6��7�d�w/�����=-�	�w�z��U�<���MQ�f���z�0�����8�N?u-8���Z5.��:���l�G��#w�Ox��%��M{*,#�/t�7�f���3��j�EA�~��!��-ž��TY/���cԎ�#�EWEX��&1%=�u[���p� ���|y�9j�Pm[�m(YA��eA���]zЫ�y��7A�%=���/=^�5V7��E����s�~���>�IS�+����&��T���W{�I�F�MK��0v�> X�Z��r����ۅ3?}�aՎ�dX>�EvE����
�#��' �*b�׳����s��`6�V�Z�uie�.�]{��`������#Z꜆(G�g]��t����Ci���Rҧ.2d��)�:��+�Mm�5�N�"�|�c�}�NxSP�>-Μ��O�q?�mXX��1.挏��bE$Lw�*�Ӌ�z繨�J�qX�A3�.�0Q�z��ҥ�hb��'djƜꨙN$���ْ���k�DRL��U���b)�y�DE���L���:<�IO���7J�ZztμMm��\�����w�,9>��&��㴂�%5���6��o�`����&�َT��sC��Zp���U��{��6��V�MM�@<N��D��y7�%��n�Z�B�m�/1��v�m��X�8T"�<�h�,Tݷ8s]�uI~�՘�½>��/�oX{��/q�m��!dQ󇥦�q�c #�o��"98��V�N���)��`W�A�8K0���w��܃������LQ��'�;��A�T�9}V��M��r^iV$��0�Zwy��P
�����UhP�I]���A��E��W�^E������+�ȡ�Pʖ��h����D�a63�N>��xѶ�Xh��ۋ��V}6�}�)=�?�	�0���$o�F�~��i �2z ��U�4��K�jv~=~������6��ʯeR)��>�Pn����!{���O�KQu��'B�X���qb�A����&A���t�
�#�̝�����ts��&h`G����j�9
<$	��2:ק�V�^�h���~G�Fp.����a�1�A��x�@K���( ���(�/m�gD2��k����f�V���I��6G�h�4d�(!HH^���Ӗ1g��9U�X2G�{�u�.�*�Ciή�Meg��Ƅ��L�aX%lR79W%iYB��W��	�7GP��C��Y���C�j�Z��m�~O>@P�_ĳؽ�	7��^�BC�n�ˤ��Ɋ���/��p�)`��_�����`]�P@�O���;�г�a�����q�1�Gt�"�޳��n�ٛ����≑%h�(K��u?B��C���ʹ]�4�0�K�{�~�]�k��L���Og�yK�������)�M~��O#vG�9��nD�'(=d}\%H���g뢫�.�w~�\`@�����i|�dt�n��R*��x��F�E��:.������s�F����SaM�*��?�U�󀋃B��p��3��rm0�����S(]���E_z�{80�d}ŭ*,�#�t�,\ ,8���a���t�������ti�S����Y~���w��(�yע$>(o&b��O՟��H\ |��[(\�B,Fx��Tu�X�%�?I��֜}M���PԏY�a!��q��,b��j�j&f��`Ɋ�S�徍���՛pzd���%6�=KFcԭT��語��mi o����$�ȱC�x�Ew�Z��AuN�ùͦ�}�/�5�hK������~�WD/��7�ҽ@�gUX�Q�$�,==n��O�V�"�Tw��d��*�מ����Y������C�YZKO�k>�^j{!�>����R)�Vj%f;=�3��Q�!��[�Uc1�0�?&O�F���Ԝ�'����S�� {$��m�0y(F���������k��PX�b
Cg���Q�Q9�WVvxꐘa��Y�v�0Z39�_G������f��dySXclJ<�7�=#UX,%4��H���k���b��?�"���S2��(�%LUF���B���G��a�<Kz1�����(u��s/�Sp�ߔ�F�2�QܚM�+h!3q�ޱ�͞� ��@߹C�*�n�w{h���d��f!E��O�
�&&r�'�:q���|�.�{�~D�V��y(E�Lv>��|!�w�V}��9W��Z�<}`��L�gx��b�b	ٲl=�¢!�񌐐"cE�<[�~�ĆΆ' gLbKxQ��W8f}׊�\��P�)�7�%/��C<0��QJ؋˥�8�� ^Y�N'��z�+��WFɖڬ7��y� bO&�XyG~�� +�1S�l��z(�V��^���t�!1�C�(GZ�1�
�W�û���I�K��`L�(�5�'�C>}�#�U�Awj!I����k��q�9}z����\�27�4���}IY٠���rN��B��ڹ�
Ů��@!����蹊}�Pd��dC�T�Oǯ�ԄK�F�O�W�����Q�Q�ŧ�0�-�[����a�_E�٧��A�[���*�r�;yŢ���b�˰��QxX�,{y�
Ag$N.'��m�'��wb-������aE�����X���'��N@��,m���:J���[H���j�Z �x�J>㬃��6Ms�mx�^q�aQ���ʢ$�ÄtZ߯�� ��~���gfH-BD�\7�`e�e/AoG��~y1�#����v�UPXʇE 2<�����Y�����'�O=���H�� @������h�ḽE���5�( ]�f��J�t�>h�B�/������9��4I��mD�B�d/):bA/����S*r�wMz>�Qz�,JZN<�`H�ݝ׭�u�p�y�op�oy���j.KO90>�I3%�`����k��a��jO��A{��)/#mw?�ֵ���W�]E�d�Z-�PG�mǪ%yVe���G0����E�æ�����bK�D��a�::�l*Y>ޛ��H>�D�b�םF�v���8&��V�-��6Rs��������4��p�G���ݎh�<>�=i��G̏��\+���6�y��m-��&g:�ǰ����ʠ_J��A;��-������1JO�m.:�;0qS�"�>ZS�t��Ǖ�Dy6��7�+w��ٱ��
�%���$8ښ��%�gUk4�%{���� ��k�1��kͿ���i����L��O{5�ץ⊠����,?=����Bu�:�Y���f���jsa6��='�@�������O*���J��+ 6��<6ى�j�^g�g���v���Ъ��_H� ����;�Xf+>�r[R���"�a'omiĀ��ɫ��&�㫾� �����o�îAv.�hǨ�A��}vr���iAN���] �+���N�a
G��^ܹwܞuA���]_�Nj*��z^��|�"��l�Vq��H�n���0�OßV�MI�s~��ߛ�&u�1�KN��$Y��I�(G_����)i�u:-i�����A�p��G�8k+a-����$��;��m%!0��h�t@�����e>��Y�ס��K��3�0�w��Ad�Z]�[u��Aρ����J}��+:��a5��P�k�$�+)E�^�K�;55`��Q4VG���K��p(y"�w���yoPH�5;Z~����.�
�Z}�qJX�Hˋ��t����%%J</�8ğ�'�5�^?��D�<L>mn��C��<v����g#q�?8�A#1���U�4������6G|�@�j��h8Yo��gyd\D/�����ࠤR�KB�srkv��w,��vw�7g�m���=�<�d?�n�%g㹺ߋ����ζY���5G���a `����03ԦT(נ�.�k;1���lb��q�)y�� �BBh�vv�lTK%�*&
��q+
Zڑ���c~���,	q{���AH��j��?=�2�E��b4�ϼ7�;�����G��MJ`%"ߟV2��?aov�:�l>iu�m�5-��P%'p��5�3y0)����w;����K�ߞ��5ptjҩƃ�IR5���B�,�JN�k�=UɾȪ��S�ACBz�$�jV�6%�"���t7��ǁ?X�9�Am��K��r�1s@�W+�P�ME�3�4��[H�R���d8�M��-\O�A��F�M�4��mR+rK��b��bP�τ�G� ��;�ĸonB����5�Pc�S>��� P�P9c���,>������W�SO�H��?v����V
C~�jY����5[Li��i�c]����&��$�F"���r �at���_}4n8�����c������8xb7��71J���dM��Q��y�Ԣ�މ����/<UA��6{D�熽�'S��d�A��Z����MKI�����i4�n�J�Wٹ���^����`�R�`�Jg`�� &Al�0�ۮB���V���g;���;�(T2�Y_�&qd��T�#�k&� p�t��R��3k/d�־�X�+T�9?�\ƞ-�Io�{c����jz��c�R/�W���Kҝ�Gd(l�c��T*�y�3�t�R}L��nDƉ�%V3����Y�ʀ��*�Ax�h���j���A�$X�T0��[너mry��5��+ ��;V|�+��o��u�W�H��w�o�2 m1*���hSK�]i�	G������s��4:N.q���<Z��	&W������a5Gۯ��D�Û���I��0zy]�#�v
Ob�c�5��L�h�0<���2rs�'I=����p��ތ�M3����=O��@m�@K�F'��ɦW}�ɗ���hY\���
�KhGdY ��V�I��aB����4y�Y��_`U��W"�y��}�.�gND�ǽ�
9J�-�z\K5�"��v��2'�Y�����G,���ICÄ�t��3p�=���dz2�I;@>� ��(�\8Q��1����J�+���� I��X��a
U��J�-E���$�7p;���ld���/^b-�������j>"�[��O�-F)�D�h�G�X�fm���.���WB"���a`�����י7h�3�)W��ƅ�5w:��[�`
���N8*�������m����z��3�� q6;��B���͏E�i�"��Q��&4p��	�z1WI�G�0�t��1�x���YO)b�ad΂d����;����A��jJ�lXW��S��V6b�Fr�T��ح'��z�^��W��9T�E Q�%@^�eT����p�Vw ���9gª�����>>�X��vg�«�2Ⱥ���Dˤ}�<���mF��:����FJFJ�����
Xۣ(k��&3HU;�3:$�5|z^T���s:�|�21�A9�z�>�M~�]��7h�O��ϐ���;�߹w�M�/���p�"Nr3%|�m?TVɍ1ko��y�Q��{A����[�
؉�s�}C-�f������+�����P��L��Y\Jcz8�򗷿m
D��2����+�Dnd.�j�����hCح|�y����#�4������;%s�#*y&j����S���P�M��y�h�Up8����6U��9�0���B���;��Vw��c"��j���Ug��x'' ����,9�9������	�`�%�*�`<����� s+$�~�ZC�F��/�!�)(�X���x˜�vCx����y7���)��Z�e�N��'�,�4gL�\���)[�&��.�QXH�����+1* R��.���zp��%_e<�h�}O��,�\h ��Y��I����%*S��Pj��zK��x/�!K8_���¥�����|�t�Q�C��I��J�%�Ԏ����3�����ʔ)
c��)�qx{�FZ�T��/��l�3\���w�&!.��������z�R��V�&n�`�����~N׌��5gw+.mQYQ<��f{y~%������mݹ7CoH��"�a�?u���#�����g[X�ٰFF�޿��E{��Uu���8��q�[K��s���lڈ/Y�M�������mM[�Ok@�*��d�˗�U�cTE�M ������^xG�VJ}��,��xÃ���z4Pj
�)8K�K�)XsGg*�3��ȝ�_*�r�yZ����Dq>���d���Zi_�c � ��q��9�9?8����eA�P��A�2MY�������k~
V�i8E4��� �r��/����/�1��y��(@ Z~����I�Biu�_�����2|;!���,�	��@��-�e3��j�B1�$n��!�oz4����F;���i:nw4����N�vů̋���n������0�!2P��s`����	#�b|��(p��4~�goI�*��NQhj(��5es�Lj��NJ�]�L������"͋�аb�Ս�uۚ�me�PQ�H��h<?�:9h6��G��HWB$���G	���UuU\t�~O�b��k�6�=~�;A���:ȰɫO�v]ե��?f>�j)"�`�����	Ne�C�E�7���u�e�:D^�Pg�B��#����m<� ���S}S�d���ْiO/�Jx�D��<[�Y	V*%�x��J�4��U��gX5n�bg�A���v�c;f����5E��f{���D�*�.�wP�u3R�|%V'��1�8��AV����:��}W�� ���?}�d��Q�J�ߜ_ձ��E�,N���x��A�=�^@k2�@��%~��B+�V��������J�t�՜	�
�C?X)Y@]0^���?�`�52��!u�O�	w���U��S����.Xg�O��RxD�g/TF��I�p���B��j%l61 S��F�&���[2r��0��*_��y6utʒ%h}+f�۪���\Tq2�������������kf����V�����;�;I��{�VX~���9�������|_�5�p�C]G��{l��%:2��`	��z}0L҃V��a��e@��m����A�y��?1}U��WR�.Zy����a{�b7��XE�3r��/ �š2����>Q{v��-J�"4.����ko�U�6��~ۛ����fn�[*��W�ݏ��e"�-馋�����q~����U���\XY��7W���Kp��[R�[k65V��%��V�6h���Ԙ-n��Q��c��SHN'ec{1\s �p^A�z�<�#(����C�.�NO������zy���l)������j3x��pD�e��A@�`>J(D�:&R}�K�Ʌ��QܓG�/mh�V-�����1*���{Yи<�d�tV���8���Z�/,���Tz����z�Y.�rS�d��G�f]�UlB�M`9�<�*E�􊲢��~�*��:�`\6��P���s	�s�b�V�z?�2�������{�)��p����9�&�� �T`$�+ۉ%�uQ������Ʊ��ƶR�Oz�$�a�'!�'))��ZmEr�s �8�#�C�$�؈�9�=�	�>�hV\3��D�u�A�Q��u8YI�$AH�+�����}�F���V�34y��U��۹��x��x��U�����)�͉\Ʋ�nnõ�d"�6���r���a��X�P��}[5x� �&�Onf�!�$,A��|s1�3!(�?��d�$,�0�q��acF��	hL���>�*�+~��e�4�K�O�_Z��$�4y���&��f��hp��(��VUJ\�v��1��굶�v��Bs��hkV-�-�:%Rl����p��������T?5=��8�4�9mό�}*qfo�iԪ��������sU��ٙAȕ֞��D�`˩��ϙ�6��	g1 8�)ꮲ�Q�;��v���ܾZ5Y����ʌo�9Ց!���v0t���e.�2H(M]��թ7�U�,�:,W�����k�; ��{�����3�aep��ѣ� ���hGe�V��|,b��>- <�D|)y�A�;�K/��T������co�v�:��2���s�1Y�U�'�Rٜ��ٗF����������j��f��p�ec~g{�h�H��fh��Je|ɩn�A;Qz}��Ϝ0��z 3�J��Z��i�nѕ�	[@���:�M����hݸH]Z2�9( �F7s��TaB�Z>��w�4��<��-9X�\&a<��v��sO��B�U�]a�-����*s4��N���*�[/�'�v� z�}�����4?-A�>B�-	E��}N	eȽ��wY,7�w����(w�침��0�`[[qH�V,q4�1�`6��N���
�w�I�Õ�B6)�XeDV"�ŭ�7o,�ſ���MMb�y�)��&�YY������Y����e�i)@��Fe�ꀶx�2���-�j=������p]��������t:=ʔ3��״��T������U�6����h�}d�[2ki�đ΀�����q	��s�4�Q|�D�
dғ*�O%���(ެy�r
�H���ֱ������m��6 �Ay�	Ur��vx[z}cT�SV����>�ζ@[v��Y�8�[�۫�^H@��L���Vt'ȿ♙��w��Ap�=�g~����!�y~�Q����́�Zeu�1��Ȯ$,����e�Y�m�T�8����N�2T�ӂ��AN�(�hg�"E��˾��+>+�3z��'Jk�}�N�oz������"��6�����j�b�o��x���Q�	(��ɠ�e�_�ൂ\m��r�n�7�Ռ8jo�aˠn�f���@�F��CV�� ���e4�@	CGn�"V�;�?Ks�Rc�V�ٻ�}M+|�����B���v�t&�O�#�>I����Z��	�62.f�}��Xd_����ıbD�@�h�����e]lj�8C�;0�x_	ƅ:�1pJ齃�l[����Y:r�?rk�]giQ��lh�ȡt	w�R�H���X��8���s�2��:��s���� ��P�f{B��TXd��bK�ގ%"��N÷�`�𫛞h��|:ql/~T(��މ����{r?�Z_y��͋8�W�-�ll'���b8�2#Y��]Nس��.ܑL
n��+gಭ��!�N)�O�죒�m�m2f�A��Jx��N#N��J%5�u@��Z�&
b0��3Ƌ>�১�L������s+
�O:Kxϝ�DU_�3�a/�@o%C�Ask����|N�C��_/�f��93 �i2]m�s��m�`X���KSI.�����?
�|���Su�9���jP��u0+�_�"lU�{���MV��z»���7�B�������K��g�pvQ�כ#��i���b-��dS�ጌ��{߶�9sI,��>��7j-\�>�yď���q�#���R�[Eձ���K��]~����(;�@�1e�������,�� ^V)b�>�3������7=�2Ӛ!����aD�Y�_F<�V��v�U���i:�geߋ(�O���JU��y�Lp�7�	/U��r���w�d����x.���3;̼�_�u�06'_S�+d�;�,_q߉w<�����T��iJ�@$"�dLpl��xkE���V~\���_t�2��W���� �.�*5���)����ߥ�񏂌2?��KХa�����b�4{�2H��^����'�;�m�@��5";�)p��]�zm���^7�wˏ�Q�AY���?����hZ�ŕ�����\I��om�(��V}���,��Kv�v�<	����H;�Y�v���Ņ�q�����UB�<��ص�*�<�� ��o}��Vuk40��,������	�h|�#�ק��Ő|���E���A�m����d2��(��|�<����� �.Pe �/"���2��'����ᄻ]G�$b�i��1Vq�h��L����S��E.�R`8V^8?N�DE�����c�1��`~Y�s�N��I�٣W>2Hʇ�.�UX��B�F|����}ۏ��@0$�и=�ؕvu�Y��F�����,��c�[�G�� �'�fM��.��>�op�X����%K�=�$�)g*�Ëa���em~����n�y��#{Y%�)0���5�:R�눣��+��˝s���L����]N��UW�w_�l�t�]�e�mA��-�I����i��q�.��1Q�p�>ˇ�-�jSS� mC�B����pMڤը7�dS�А_E\K�H�������q�9^���6)�6��?�(�!�DئM��Ê��H�}�� �sH,�Oز�7�_���F����0�\�D�LyCE��%��g���*$m�S��Vl=������k���pB�aӊ�g9���<``�����M�<%=�-�.L.G��N�@��ڪa�fh�<n��Aݤ�cĭ�M8d�8F����L>�9�j��aب�>S�B+J���2�����M@˷5r^���ⳋ����Ό��[v�E����U:���6������|?lA��]8i��&�����@;��'��Fr����{&x<Em+L���4ix�,`S&V�Ǆ0���s˙�+3�"J��W^�N	Y���'�hz<~㏪6������e'u!W^�J>�Q��n�Ѝ[����]�	t쩻Ĝ��W��!��}v��b[,�B�ޥ��R�̩Q���-���v�����K5��}0���~IO��&u�q�lꀻ�e~�4���T���fApY��S���k���5h�����<ޢ�v��?M�b��B��ڇ��n�7͋�O��q����9@���QF�����K6��,Y��w{����KH�� �}��ʤ���[-� �������0������]|��vU �J��oY<_@��!�]��M�4c|�
}
�e�m]���?`�����b��N��rq�%J=���Jl��%��Ru��F:����H�Q�K��
F'?���ﰟ�^p໒Wy:���,7�W����2��"�*�
ea�N�at�J�W�G����ɥ ���b�WU��1e(9�o?/�-ڇob��*f(5Tv��x9�Lٯ��F�ӷO�-����t����: ��biEP��,����~�&Q�๺g}����%�����\�nU,C�5�g��(l)�c<w�[���Q�
��)]���d�N�[��\*�0��d(1��d;Q�/`��qo��4ń�:!��2�aR�����w	K����	�4о�TGU����֞��-
o.=��p���
[=�W��%�(ʫ�C[,��B{����%�J��O�bK�S��ZԬ{9<aV��#T2�kJ�m�gFhd�9�F�\�l\������Z1�/hެ��*�$�2g������%JЋ��X%6�3I���a��x�g���f_�۱���ֱ0�l��V	:�D��� �Y�����&	m�g�� V�sGS�~��߄us�9�$�V�:o�ل���INQ'�qBYZ�<�4�����DC��w����CI���5��'���m[8dsk���ޕ��ٺ�L�6�u�մn{@���@�(8Aƅ#3Df�'�BqT��(U�5]vP���vl�)���v�t�^[F>4J]�X��88;�|�T{$G��220�����SC�)�c�h3�/���y6��*{δ��G�����/-�a]Y|�b �S�o��W���P�A����ϝ<���Ə��L��)}��-��������M�*J�U��(�˷T����=�Y)'Q�L�Y�*ie���J6�x�X����@}�^zZ��	B�P������
~-�[�`����|_�,��M�ڦ�$��1B�;��K>1��1�I���_ħ}�����0(J��T �vy�X�gGP�$���A�ÆU���S�K]0߃�(|C�-�iDmUa���Й�End����+��2���=�.:K�w��yL�y!h��IW��F�`����QW�Q~#�Vt�;�C�Gj��ZM]9��~�	��T�>'ջ�w��,���sܐ�x�`"T�YHQ�E��.�β�̧�TD\�L�Q�v�ː �}��N��g������NksYU67�D��s���S�5�P�JD�T��.�d�7��V�Ӳ>��pA�M �keX�����s��s3�j
�Z�^zyDM�G���1XK�v��V��U�"�'y�l��Jz�H<�B�S�����R�5�����]hjV�S��J�V=/��8��S_�F�W4�$�0R������/�����`4,s6}MG�s����brk��|
�D	�6c��!��R���?{�=~THH�O'(����T	'�q�ѳ�t��h�%b�vig36�ͺ&���q�E�4��z�`��^��8��'���g��G9m�6��+vP";�Q`0���m���@�(��9ߣ
��7]����'9�Rs5E����Qȩ�B#��Jy���c�OX���ؕ���V��qk�S'��w���6��jI�SS��,�?�������6�|/ʞ.�	�u���U�����-W��S��9�St�}7��3X�>	�9��c��9���2L�Oe�y���������#?Y�=)	m=��Ȣ��3;����Uo�Zd����FG��9�$��T1iD�lʴ��%'T�2V)��������&8e�^�M��W� ��3' ����e)��������p{o�8��a\�U蹱�f�~���u�([o�yT�}NE���((���C�`
]�����ȴ�_憏�##@J�&;D��vBƻ<��LLuz��P�+=�
LN)	^�-�#h�>�� ���wm	�V�v���펀�����FAɋ1��N�14+�te-r��ͥ:Me!���p�A�ץ�x���>0%g��n���!�N'18'2����y�=@��-�i�Y*~��ض�i�>Bsa�$�*���u��g��½,��q&EI.>��Cb���絉���������to2��KX��F�b�_���hƭ��ix��l�h��r}T+�3��UKy�?�f�*u�]=
�9�y���H{$��b��"i�5��|1���ʢ�J������5�خ�x��aڥ�|��ƨ�G�k2O��cA����>0�:i`����`�\�R#K�����<��BZ`�%�q
��JؿG!k� �����YzKx���~DY�B����6�rr=�� p̈V�6у���+㏖8�
2%�?� cdg��Z����-)!���� ��x��J��W���|��F9f����48�E�'�Q��\�5�q�/7��by�]P�2�A䄅:� ߯�� 7(�]�,��CF��,^Lc��
����Ä��z@_��@v"�b�ᇺ}��)G�M�#w(E��JF�-g^�ݘ���:șP ���7�eX Ke$��7�%��f�"�?K��&�$[�H�	#�24�K0���o<��Y��6�,�E���MB�ж�M�B�ti�ym������+�����rx]Tx����S����:�`q�m2<�r��H�2��^D�]K������>������tיc_`o�`y��VȽ�Q�4�rȁ-��b!φg�:���Gb~|�eO�Z\7i��xcD�A����K
,=~��lND�җ)�m(��+�JI�=���a��Lr�s�r�"&΃���2�� ��hJr
�W��f=%.@o�EV���H�
���"텾ӋmA�����,�F1w^�!T���0u�"��:$�TKe��&�̴�y��� �w���E�G��-�;�i�9���v�nv�
�uH���_|#�%n:`6�����ڪ �
 c�
3�<���ī���4PG�IN�����RS!��9Yk����3'> W^���,@-�.>(m��y��?�X�Ns����a=`�5kT+�[��*an��Q���c'��dж�|��^��n_e��)�Cɋ��'�a� ڹd�V-�3�LZ!Ɓ�0Z4���@�єJ:�c�f�$�z9�K�e=zu]/4P '���f�0T��	�;�/}�,Q���QQ�;R�����L���YGZ�Hɜ�����iiIjV<k��|�p�g�z���~@��QM����

��ݖdp����z���=]ar���ѯ�]}�a�6��v�-Y����S�If����A���j������)��!�Քy������3�{�1̥"3�ƍ�jPe&��}���"u<Bƹ��E=��zW+�(D������́ڹP�r�I��$���Mm�*J�s
[%++�� ��s��EN�Kѡ�(�>�\��^.��W���N�X؟B�,p�'��qs7����1�.:�{F��lg�{' g0�S#X�./C�;̣���I�c�Va����EY))1�m"[�l�,IG�
�_T����d��{B�i]���8��1�2�82i���6��k������/��J�ՉP:�O���*�NG��w�|r��@i��f��A�Yw
�?�7����z�R0e�pPk�4�������\P��d*Ct`,s�O�-sȏDI��g��c��"H�\9~;������S�/���qq���č�'�<�(P�E�!��I������Y��|b"�?�#z������2���>g�	M��_>X�;BZ!�@:-�&-�UlQ�n�A�ä���_!Zh&A�p��O�����?�b��(�Q�I����_�,�����.��r�&	�v�g�A���E�&Lq�bK��=�j��&'y8J���zq���Ae�%���:�t �#c�M��Ҡ�0(��0(�U�\���c_"hK[o������97���,)�
�!#Ѹ�Ó��d;m֩���?wO.�(+�X�brB���B���x�g������7/�����j�ӻH�A?�I4!�*�-�@�	f(N\�����H�!Z)��ȯ��ᇙ�i�����
�~�����S<{*��8����$�j��zF#z(����q�[������ ���q��1o A v]M�bA�����q��q�m.�?�0��7=f�tt3w�1\rZ�uG3�u��%�1���`Z����|A��J76�(�~=�t��U�N}.�ȇ�*��{
����$�Q=�ɱ/i~͓̊x/̔���2�Wc����O��Q�'��+�@�Xm��dn�XK;�~�H�&{�/
E�9(!�7���< �2���5Q�9��P���s�E��qn����T�'l�2l�lJ�*�}�A�x���Fā/݋ܽ��݂?^�oh:Jե3�V^��|��d�5*�j<�%g�dp>.�*��4�^����� �����M\��^����7�C�Y/Dx���㊉|
���]@65X!�-J��ƫ%cˍ��;��K��RJ=3x����p�oo���1����N��WV�J��!�D_���]5�#?G6�1�;���{uOzY*ATxYY��=.xh5~켻�ۜ)�.4�Bm�����%��2t[��� �%���I���zo�5���������u�\�^d� ���u��ϒ�r>s��s�L���\Mn��s�+���~����<���`|GH�4b�㎞�����'2iS7xT]�M�)�5<�2�jc�R�N^[PDCT�{��u]�<�N�f�Y#!=�ɨ���a�l]C�oa��>�8����G$�zͅс���,(��وA�Ir̈%E ���^c|:a�gk�rS�Gh�d��Z�<PG;�QH�΅9nU7[��'Ӓl�xZCԤ��cV��L����o5̙Lw˼%��I��nOH�E�o�V�� ��UMҶz=^�؞I�q��ZO_�tF�Q�?��c]���#���<�W�4��:a=�B��H[��`8����0� m����6f�h�L)�h���۶T������축[��2\B^��Z��D�$B��L�>o{v����2�挏(�(�ɝ�C�v�6����ò�EJW}�83�2&����H�ʽ�+U�u�є�k��X��EI������K��@�8���������7r`�D�y|S`�o'Wl��G?��oj ��M󉈲��Gt���_��+՛<�촩��e�#t�y��)�����3A��c���U����4N_�D8��uk A~�v��@%�jʛ-Z#=�������fg���CMRC�����fs�
 cM>�;��MŔi(�x:RVZ�1a����E��
PL^G�N^@+�A��~�g�	Q�e�9�Gco���C���+�������F�ȿ�HHx���E�x?�M�I?!U�C�rk�7�㝯Lٰ��DG�)��LE+����8�CU��x�%�XӘ��u$t��l�P�M�Fb���׮_��$aj�Y���t����k���׏��U.//���V2j\�J�c���<��x�r}~o@��N��j��	?��S�����ӇM�C�B�1TYT7_ɋ����Q��9����\�J����/3��z$I����{H����v��[�%�>l#���m�/W����[�W���<��.}66���^��T
���Օ�2س,��R���J�I�N��bh�8��f�6�X�o�c5ϊ�Y�L� �ҕ�3b:��妙vX��o�i�Fʯ||�A��O�RC����@�[�F�-dBB�
Ù/�� =N�f*<t<
>L9���i�}����ګ��S�21} ���lO'��(m�M�J8��ԟ@�p�e]�xq�\��?1��,!�_=H��5�YO��.b����;O�ano��CpIaOH��3��0`L�𿀠\oEz� ���+�|���==�@wf���-��;��f����̖��x�;Yau�7��p�~P �ݧ�hw�4/N��;cD{�a��m(M���*��̫�.;��;SӚv?��=�}���Y8��@�],w��D�F�yc[���`k`0�����Q���4�$2c�3�;��Z���96��vM�!�agPA�a/���!����E�GPL%�=3���/Y��}.� s��Q��5-�F���B Q�B�;H!%F�v '9�2�r}�M�eW֧w.��$ZI�|�#R�:g�.$>c�4B~���e;����� � ��!U)���_��H��,L���G�e�0(X��)���~�*�C���⯊)w�'E���u.E�#���b�,+D�6�Nn���Q;���� �)����Go
;�[vi�_H|[T����!�s�ހ%�BIx�k�N̞�}��0m[7>\�7%f{"c�";�Cd[���4{o�7yж��Xɂ��w�0: �<�O���1�9��~[0�
�����.�_�� @[��F�^&�����L}��J�o��ܣ���,*�\5Qh�x�y��;�w��H���:qF������E$�P�<2L�%ٻ����F�	��t�Ydo��3�#�]����>��e^��x~��l�E�Wx�9@�Ѹ^#aS��	O�=��9��p�E����7e��7��f%��[�0��q�.��B�+)3�4�	�x&����ֽjpͦ�$���_o :��!���Y�^�R[y�X��Pa�p��
�8D��fW]ls
H�����/!]�)��*aX�2�=[-vW{1��DG�~]�������nn�[��kE`i�TX7h�����$mF�ua.ՓPEG^�R/z��~<A��z���˴k�J��~K~E�b��^q��KOQ��f;��./��R�c������yv����@[;�%��:"[�!Њ_�
�v3��C��-u�.|?�.ǋ���sk�j�`m-`"!������?é̙*$`%��¤��|�)���H�W����Ȉ�<1�"��r�w���
A�"� �ŴX��?֒��8��>����#%W�_#�����ֺ����*����k ��&�O��:Ϡښ 2ݹ��ə�69�h���ı��(w��U�=%�<�����jn��VZ^�	�qȋYKjU�r�3H�Y�����!�g!����B
/�}�Jf�[�5��T!<#-�z၍)$�aEB��v�8y}�\�&�����F��X|��V?���:�W^�B���i?���%Fd҄�����u���}_d�Q��"6�ʷ=̬T�t`&{!��7����,K����Cgax."G"f��~o��Ƣ�]��A��g��Y=��x|v]����Շ�i��$��HG �+%*MR���)K�*�����g�؈s�P!K���	q�[Nw��6�K ��}*L�nk?k�C6��t&���zf�ϓZ���ۥ���Y׎�Jd`P�9Qpg�/[�͍L���&J����A���]��t`@e�LW�����k@�ҭ�	��Uڬ�c芵Ҁ;>z�'I��z��{�TƈnD�b�"��P����c�7rh���ыZD������|�i�E����j���mgr�ʆJ,%��3�^�=�� �j���ԯJ_(+Bq�$t��Х����S�� q=�˪7�y:&[v���؜-b�є>���-k�SA������̑�h�N�җ�\�%�7����/w)=}�jWY;��Y�	�0�+=q��Ð����ZK��ѕ򲓇��g�B_=Z96�u�
< &�c=<p
�!d|JC�G���̡7��Z�ſ��'-a��g��?9�i��p���J�l���E�)�h�����f^!A�NY@� �Ax�p�U��M��?����t�5��������I����-B[�[ꀯ�l��%���*��ߜP�]u��p@�N��wl;���t2rέu�%	�"~���{�l&cP=|k��b�EwW	c\���n�n K��ql~f�&L+/�8��~1$�p*�oj
���tR.�G�_�1��a� $T���a�ߐ��0�����p�����齈"�p��q�l�%�ss�hc��h'$,��	�K-�&ˎ�:���.�>d9�a	Tt�Si~̤7n���ֵ��$��3�
q>`�"03�d�1�Yz�[Ϣ6�3���&�CJ^!\6H@1�����!+���Z2!6]���O���jG	6Ca�r�՞�\�R�H~��$��"�V'F�Sf���ʠʊ��I֌��s~k9A�q�^gA5&�`i>+���[���H�}As�'M��Oţc�V49&h=R�V�O�ƶ�
�2���q/�w*����Y8�lҸyg(�W=�M͊����ϳ�2`��\��Z��/���5N�ԲD6�gv]�+CM^ԟ��r	�0��k\\�y�J�f,�	A�}�MSY��B�n��d�J��
�3�a���Bv�T�N�g���)0��h/�s�1>{%��������f��)O)���u�ۯy,Gt��L`�'�&�l0@H붇4�馐��u�x�H۞y�kө	�� �V�� �uby�	� "�C���zOL��ۆ�>8$�a{Ԁ���\��i~�S�V	eo���U�:o�k)�u��+�~�d��!9ok([�"x���##�.�4'�=�IT��M�o�| �f;��a�����s���7F�
C�?����ݱ,K��XXe@V��Ԩ����N}
��������fS�~J��c�5���&��hsj���Z혳����Ӎ>S��z\�����; ��xQ�[%�~�~蜰��o]r�J�%��A���	�$J�m9GcQ�4Ր��I�J�5 1��`vN����d�(���k;�Lm�Q4�� �C\�Ytu�V�AWw��IY>�"�թ����!�C����AS���+F�k
(��S�����2�w����j�"�� �e2���]<���m:4�؇�(ʺV��a��:�.2�����*ƙ�O����{&5�e6���z�u����R>l۲eq��{H�^:��|���#�k��4I4����I��ʤv��A*�RRw������aY�`TJu\a��FJ�5O��xgˎ%��q�CxLwa���LY�P�c�" ��cw9�w�����f�-_�`�.}Կ�SF��Ճ^��Uɲy���(^�,1���Obj��6�2n^"c�
��ucQ���^��4�zv�B����I��K �AkQK�"�Y��l��*C֫À�j�3e��DG�p�匟@����*�mI�\"Y�������¡[��I���z"��Y:=�1�meD����hh=ˡp�	z���Q�����f���n�����4����b��*���S��i���lwH\�	Gb@Q"�u�g��$��S�Sx�KyeLt������PT������N�ب|�R�q�Y�>+�[�fGz{*����tl��͖�M�%\� /VI�k����|%�k1!��i��G�v��xn���,�� �05����3!+S���Մ1��7ߖ�Ex1d����]K�����0ˋ�b����a!X�/�wt#q�Yٛ^i�st���\�?�2`!xzuݯ����/�3i8&ѝB�Z�k�4c���?�c�J߿���\0V��?Q;�x�h9��m���8J���/�P�e8|>�erH��3�{gxU���t0�i�u�(�Qt;(�%��<�\J�i(�����r. �'}�Cb�J�7�i�9REXn�d���c�MjfZr����8���s5���r�	؇���ECg�Ԛ/��d����r"L�3,Nv%1hfΞfn=g��w�z?3������׈Ͽ)�0��HYi�(���ؾH��?��+�i�7o�<U�[$�-v�+T����G�����ȝ�H6NI��:�C�Ϙ���tŉ��Kq�d���?�1[Gb���gY&�u��M����V�|١�IE�hư[bA��M=��_�u�ML^�������|(J��aPܱ�C�\�s��1�Hnb��ޱO��=�B�p�����(�	3'ø7E����,�YB�_��I�:^�-��&\#�z�2�lLt��6ֵ���h	�WUm�֪n������=dn�Jڤz�ש#�D���m��t�y�+��B[ɑ��g�C����082�y��n�ϕ�P�s5��3߁�yļz�>g$���ٴ�����??������_�3�39��=�QS�G�){pM*ƼuvH(?� K�.�w����msq~�V#5jwG���|�aJ�y;G�[������VQ���/_A��2��	I�WKF�^���䈙qF�o�	�{W�ȸN���D4�� 3�� V���.j�-�$R?�5���DmQo���J��/�n����'�P�k�ԥt�t��X%_m��r<�["��0xO8�ëB�^s\����C�	Be�C!r���厝Q|E��w����P���"�%\�O
a-U��	���dES+�+�o����r�F�Xآ�?�>~E��W�ν?�7�����&�d���8I��^~��~!l�$��vt��^�%�v��c���U���2'���\9f����1`S��]6�(l`}��q�t<��Q7H��8�)��q�H:Y��x�dɋ[�:�cH�}����/릶N6z��MP�(�p&��l��u��8�jt	��?-*9Z��ٱ����g�λ>�4�j6v�L� c�P^5h'�Lak�<̚�Z����y���!��ʬ8Nh��
��s�ت�敝βg���̣�x�^� 3����hA����cD�6%�c�/`7H�m�nHzo�t,��ͺ�άפtk?�1�	��Z��I#���E�*�M����Q�Acu�Q�4��g?4
^�D.���̟Q�dmG��P���L���C�)�1$2� KS��`6�j�qX6�4gª���xc對%�˙��d�"�6p�Y$w����xV�ڼ���_$lJf�U[v��{����?�}hS�9��(�_������&��ysUN��w��q�@��s��ĺ��E)$2�J�q�w����sO����Ύ0�y��T��G�jwfw�S�el$PRc7���� 6�!�,�r�d��P�<��U[/_g=(���M��q��-�">h橫���NL>��"���mɞ3N f��:�z��L�%�ի+�j��V������O⇔���̻����F͈2E��(y;�<�k�<�){.�)�<̅�آp��(�L�OW�D�vU�p�y��i7$�ڥ~�; ��d�������?h�py��0ٔ�#t���^衎�_�V9����^�QyHgv5X����=Ć��oaN�W��Ә��!� ;
ݤw����VL�7��Kx�dC�
Q�%�U�2��t�`��;6��=h���Ҹ&��&����I�7~���༆��npm�����H�ŀ��3��2W7,��P��zT͆|��;��Y��5��5�ؤ�:�� �xإ����~�i���k������[?0�t��|ޖ����T��[��헼/��a�|?�|#��X���B�[Cm����l�����.��wZ?�/����:7?�k��?��e'�����.,b�E����Uc�"Ḋs-ζ���'Ȩ��?V�4ܓk� 7ƭ�C䙏�B��/��͹Rii���(\�����-��!�p�0=��������m����5q�<�eKc�uֆ���b���z�(�"���,W���n�M1��Q��*'�G��E=i�69p�翣��ƙ)T^G(�H̰�e�<Z� ���Da�e犸S��!���8�Z�����>�akp�r�5c>�4���=q�R�h�<�U�9��j�C�f��f1��\-}�	%����0�MO���;p�\p����`Ɩ�~�II��"A�}Ǹ���oAHw͑�>���A{)�(�9��� �	ul�R|j�L�|��y�V�H���_�x�TdK.��R��QƩkl"Y326`u��m���Orת�����:"�wMr($wqZ�s-bI�(��sш�t� �/l���s��Z��P�`A����J[g�	Q�Vn>��$�S��.ɪK������X��;�S m��v����v�wuAv��ao��JƑ�J�pF�녺8���U�xU�G�Q?[���2L��ڜg�}�p����?���<1�=(CÜL��!;�]���VA�������0He����%���q�����qu��\΅-$d<�ݦ�{[�9�%�"g�p��b.�=������5u?6�~�ǭ�GB2�<� Q(A�Ь42��7��g��h�w�~f��B���y�5�	��ੁ��5����Xخ�r9=?)ԉ�0i��h�1�{ht�*�:p‟h$Q�[�Ư��Vp,JJ6-���lD>]F�'~���M�����EOⳍ�	�M�lf�r�V�k�-�tM������Hj&)1�����ԫy�T28+E7�lr�&�mo��	|ޜ��,����g��
/�		���ߧ3��2�:O���ݸ��K$�����I+hlô1�-�|x����iM��-�I:ݲ`�3Q�Ê�f�\�L%��(����7Gw̵-�!�*#����)ͨ�"O�l�@v���V_X%��(�|��5��5��T~�pb��(�Yq���7�dk�Y�����{���t�O���(1���?K��p�< &��C�G��Zg�c���\���D�DL���Ř�F�ф���zy��/b�}H,�w#jaV�ڕ$�9ڢ6����[e��z�w�̲��������q\��+y]|=8��j[�o���f�lI�u�+���|*��ǽ�s��W|��&����D�?؇i��}��X��D�-�6�����{�6CV���'�RE���d�MsϹ���
,5���^�h��)F�G�
#w��!�o*��~S�u�_$2�F�VC�~%�Uu%��/$�=��lP�Չ�� �x�U�:X�7��6�F/&�Fc�ѧ��Φ��=;�>Fx�)�	�j&�=g1��v��(���� 8���=�K#G {Mt(���ߌݾ��A����<��;���I�2��f�Vl͢�8�	�R4�q�1�ߛ>���֭[ւ��k�r����`�A%��U��1�U��1�9Wp�N���L�P%jV���6�)c��
��xx��u=����l����weS���r ����b�a1�mg;�G�Z&<���%u+عi��DLC���[j�������/�N�V�"�=w�9�Y�L��݁pyc�c�ڵy%�,�� Ѕ!�Q��ӣ�^` �'�X�
U�T[���oq~�Qr�,��?g��k��}~_�bb5_�uۣ��N��U���cn��*sw޿DSJ6Af�`ʥ�x����(�a3�9�����ba�`P��l��Π��Ʊ���a� X����[��"Qs�'�lL�^��f���D?g���"J�����SJ�|Um\���>ھ�/(�G�Է�aς2~��!�����p��4[|���+Cӷ¢#8�\7oMK���\������6�f�BS_dʵ�@;�lZ&5��������Kg�P�D�\n��b����b���\]L���XB�[�C_���\E%�ܷ�(;U7�o_�y�5R��Q�wäv@G?�J�!��8�ǩFƤh���I�k�mOl����a~>���f���k��'p��E+��T��t���T����7QgL�BB�]2��?���Yl/��^f5ٲ2=8�BVl�m<
Q�M�%7��������|,��~�0�Ӡ�K�tQ�ƹ`?�����$�h���?��bu09�$�9·F�6���e`�u�L�`���[�ה:S�6�,Q"a`��Y�`<ǂ���1��I0�WrMCѵWbC�m�e�B��6�mP�x4
kD���lH��uPe@�#}���-ި�^���UƯj9#�	.�����Mq	pX������LP�J��$�D-�Paj3l�g��B+���ȸ3(Ɯ�����%SE���79ɳ���up�,Y�:�����Y�R�`^oÖj�RhL�JS[" �\.
-���11�w����;6(9V�VK�����ޮ�*��d����g��VF���k�{""vR��A���R/�A���ǯ�^v-�/5(��X�^J�_/�O����3{�)�N�u��*/op���LjT?8Xa/6 cf�f�������7b�A$�l�u��"�!Sq�e -���ɖ~�yzx��_(��.%��2H���7���S9r��~��{&�``��ڎ0/c.�\��  ����u� �	�����l�FLn�����p������,�?8H��e5l?=*�E�^�=�q[=�p��
gh�_��9b��H�r@P�8��7�.�>P�w��Ψ�)�dZ&9z�r�nh�lF�O���=>�]��4���w�M�������gxx����*���H�Y�-&:o&~/O��L������S���z`���QO ��z�ռT�F��]�>�G(&u�����J3��R�_Ng<ٷ�Nu>o�!��HQTw���p� S$5K�D�g	5��A�؏�s��q���J=�$��8�����s����#���5�g�Z�,bV�Yr�`�R^���5�|�e��_*_[�y�g�j���)I��ԻZ���BL���C�&�Ҥv��RHD���{�}�c�;|Ͳ}�b��,IF�MS�@;p�%~Z����cl���X7�4GJ^��>.���pJ�k�W`a�4a3:88�	F�Ú�i���ct����>H��%0��3 2���/���\�W�uvd�I�8G�����3H��%��Č�̏ۼ,�驶�PK���$s�QsP��?Q��,@�nb����=�y�tk�̖O�7ȑ����M���/�f~���3������~���uB!�8l19�,�1/'mr���4a�]����i*k��d\�6��XK�b~�����ߵ9��{�1�H)׉��Fkb	8��2l[��Ϯ��S�(yKpu2le�K��b?�AfD[t��Y �1Z���f��J���U_�>�)�s�fA�?<�Q#��+�p?��f�(j��{�a�� %��ʩ���
�Y LH����y�]+K��D���&�.�S��p�71v�k��/�c�-���PP��@L��m��<̼�v&�1/����?0!�xX��W��h��C���I�aWb�A݀��q�m%Zt��/DD��:�\;II�  �}�v��_^��F[�8�)M�u��)`<� ��n��lr=�����H�ש�k"�Ye�k-���I"K�d�p�!��7"'e�����������@Ƶ� ��o�9��,�ހ����V�ql�_L���<��d��
�������ϱ����"���4x���"8�#��t�Cz+9��n���=
%+[vL��Y��J�=(���⣵^P��j�&R�c����5{���?%�# 
�����1o�Ǧ*Ϻ��)�H�m����&�)>C6����~!ݨ�Z��?���N8:h_C��id2<�J-��%��W�$0�-�(X6^3�������jO}*%�N�~��@��1O�V���%D3�of�΍(�[fE��4$ռ%.��?\�U�>f����-�SH��*a���)ޠ�9�Nh8^`*�3h�c��=���g�&�ŷeY��J���'���\��Tܫ�J��G�T��P�l՞E�򵇿ݱ� ٕab5�-�6��w�܅G����}�s�A1�G=���7��G?/6��z/A;B��[T슋������gu8}���I)���}_�Su�j����z�X�T+��4���`���8BE:G�?sK��l
R��_�m��������,,NA��:���:�D����k1������xW��na�yutOis�Q�JRF����r8�ϴ�N��I4:t�0��i�G�oO3��O|����d�\�t]�R���-���F�|c.���R�����¡'6%z�$�}k�e�,�P���>�U,Ȓ󰣪<v��(c�Fl-����a�B�q�֗�]�f=Il�`�
{E�aCA�%֘ʽ�?��E���QIࠆ͇|�����Eۉ����D�3w����	bԛnܣ���ձ�1�>-�%���ϐ��a����s��So�}ZE��>>�K��X?l+w�6�2d:_��E'�CJ��%�C%��3�m����US�j���@`31ڷN�m���i����f��AP�YO�^/�gpJ���c�8kw�>9Z;�ǜ�8T@��)J<���=7	k�b��[�.�2�z���E[�XÉ�:O�G�K]ѓ�[�*�F$H�m)L/���⃭�����Χ����ZU��
-IxΞH1,����-*T����ҽ��:��qL,�-� �~n-����)Gy��&\�:KL�8$Tn9M
��w5�Z�©l�}�ɔ��P;XQ��e~Ds0�|=F��"񄂭MY�B��H��������� ��c�s�Z��s��a�@�F�~�(,�2�W*���_������W)�-�����(;�F�u�܍3�Y�-"���\��V-0�#I�C�/�"`G!Tl�7��)+�K���H.Oc!/�Ѵ`r����{�v�3�E��s�
ś��e�Z_?�W��N�;�1�P�ܨ]�7U�6ne��0�\�#��.Q�#9X�5���nQ�?�t�Q�	�	Q�f=N�Y�����j�o�E������G(�L� �/C�>λ�@��,�nF�2�Ka�"H���\,�"""!��a �I��kY��.6Dp52gm��*�*ލ�r���b�^���)*R��b�;��k�Hv���;??ؤQ���L7p��)��Z`a*:-�b���۵�U$
�SYx�v�����q��+]�&�P!���ߚM�|(��Ù�l��4D<ٿ�HÈ��m
�gEW_���Z�\���ئI1@��?@�����(�Y�B��ϐ�-;C#�+�b̖�װ�Ԉ�j6�"�T��ʴ7�8����!�z�������LE�?�a-�Θx�L���ԥ��_m�0�:)��xo�E�.KH��v�b�U�=q]�ya$zQk"N*9��:�F7cA�y�VK�^�ͪI�򬚐��C�"3l� $Yf/��������ª�k����9��'$>RsRO�B�W�9�m"��Q����c�4avt(��#�{�����6*�d2���ܥ��� ���Lg�iJW�P�%Vm����b Φy���˂N��1Pl���Ep'����{v"$Rې�~��]�����Y9T�c,��h���i|���D���N�2���>
犥�4�"��h���� ��uV-Йcnxy�U��b���%
�~��O�{�������4������i���JA˛_�r�f܂\t  ��,Ē���⿾V�����:o�)Ԅ�{��� �H���~�E�:���q D��t?�l�nr�x�`L��N+��ˬ�U��et���:�joD��-w�?������q�[�W���Bf^\Q��
3��!���1���d���(����H}�H��Ĥ��m���e�NG��,�n��/����8�Tb���4�d��I�~�?g�Sq ������l��<߹�,./�
��L��V��M���L�\tG(��M��,��J�u_"��aS��a��OU때j��͗���p�M����Sl C~jӐ�Z��L{�������Ҡ���`k9dl�YN��eN6'=B-ףּ���9!�X��P��ע��DK$��i�F�n��j9��
W�C�����'�Ŋ�go�cV��ӎ��:�V����Ps�#�HYm�X���|Q�t\ӡ�P���9��h�mğ��|�[h�τ]�1N	��:����|�cY����<:��d��#������g*�i~��ۀ���� DTaѵ����>~[!.�����-[?u�k�z�\3����&���[�;@v�O��8ս%�m��{3�)pVآ�L�p�"��=��<�~�,� f"�O�ct�^�������r=D�4�\m^�:^}	���z~c [�#?��x-�}�P�j�..��!G�GSAC��B)��vAK�m�t��ۻAב8���tt�J"W�C7�ňtZ���� +v����@):A���
c`=���O���3h<�__F��O�	G�1�슦5��k_fx��X�E���̾���}��n+����h�.Ìj@�?��TlN��}rC	�P]E�R����]��rsu&x���J�é@0���X_X�ydWp�V���ВHA;ё�E�$>cSf�2�Cs�Wzv��M~�$#HZ��][jWwSW���"���]�N�/�7�'�D���Z�ip��¸S���H��}%���.�ӈ@A�獜�0~�J%�i��>Y��x��q�r~���N��*��(A�j�QYj_�8�-w�/�CbB�N���.k/��>?"@���^n��nr 1е�TU�鴣qԥ[�ΚHN�N.�R�H�j�d�
�S��e6����"8�e?&7�����ı7)� �0�`|���E.��ңV2I�L���z�$M����~�
���5�qH����ʭ��Ѓ��]��{y�ߙd�l؍s�p�Kjci,�m��|ʺ��a��\ v+6��G�=�>`���L�ϋ�4�6͌�CB�u4��.NO
�	Tg�\�����Pܩ���=q�Pas/����I�'q�!;~�'����|?,-f��T_ğ8�\�%�ج`.���uܗ��`�������X����ݮ�D��0)ލ�D��l��hY_��'싶N���՘/�p�'�v`��2�Ͷu/�&���𴍽����qy*]����HPƪ|'�µ>i���1�(-���;����Y]w�F�k/�VŞ��6�b��õe0Ύ/�rJ
�D�CvDT~V�$�w������^���am��H�Bc����2["�i{T;�[H���h��
|��ug���2�q�r�����#�NMT3���
$�����R�]^Dȩ��Gi=�S��(p�ʔ�(�.a]����8��V,�0��}����z��k\$��y*mБN��Z����}�,H�R�ݔ�y4+:|�Z���͏ߡ�"~��+�d~�f.E�]�۷��~�#��{�$`s��Ym�n��`�p`!ߛt�W1�;��~������`_��m���#�1�
z�A@F�5�6��Ɖ'��>m5�1Z@� Oܣ�7�8���$�,uE5l9C�4'چE��e�w�\?���c����2�S!�/�3�8U���H����i��	�w
Ŭ�Q m�i�����ʖ��9o�O}J�.Y�8��yQ��.����!���LK�7�/�V���#�j[��Ă%[zU�Q{B��Z.�׍S�z���]�
��s�CF$��
�p|�%��R��˴!3!�/���	}���h$	k�,`)�od���#v�\�p���N���Y�u��?@:-_/UZE�wKVF���XzAɝI�T:;K�� T��ě�oN?��F2�����.]��M6M93E�J�D�..Q|�sS�݀�F�*\���J�P:3���"y��D�斉xA�ƹzf6\m���KT1e���mu�'%�o�[nڵ>�g���P,��d8�&��mer��+���vԫw�gǡ��L���3<_�\�I�QO\��g9��3r��� 0�.��}���R[�}�6~25'�#�)#��s��4�F���Y��]t�x/e|��W����tތ���Z�]�3Q>T�� a8�휂�D|\����/�]�֫���wÏ� �I�{�ѐ;i�P���$��j%�>˟��N��@����J�6:�4T�)���-��e�[�h��>�Xz�rGA�z�fp���ؤSGM�6��$X"�I��`d_r��{#��(�d;d��O��Q��T���5@xB�>+��sd��Z�T�Ù�3;��$��$���2�%t�\w^�k'� ,��`T�h['�kl��EL� Y�r��,$�F�z-vK�����a^n���%J��'%ʉ"������1u�<���������R�։��j��
F�"��1�z��cpy�R�m ��ů��؟�Ja┬�.��D�E/IEݮ�nr��2�A�m���:�^[�CA"��V�I+Xu�-����q�>�Bv��&�@N-��	�%��"� ��*B��0.x�ܓE�3�n��?�6:�Q���i1��7�����e�N1t?�0թ���C*��=+���j�93�3�3]*�l ���i�:�c���~M�D-Y9�����J"5Fܭ�u��a2TTIE��*7\�q�F�~ @��D7���-�8���>x�d��\�5u}�� ꜯ�zGJAf�Wb�5D�$��%�t���_б�5��ӄN��;���Ġ2��IN����~��,��hCC��<N�U����JjN^SE8� ��]�5�8�V_ `q%�qF#|�1���J�T�o��$��7^��=��3���?�^�g,�4�$�*{�r8l���Q�ș�4k�QѾ�
3y__���%��=��kiϕ��#)��V`�nUW�����7+�ѷ�\R��ڜ�l�N7�~���WJ�;�;���i�S�v�q���k˙Bב�:s1|�|R���S6�&Қ��k,�Zw������t4(�C#����7~�;��D��0w�O�]����A2�&&�5RsCEe�BA�a��lm���'N[�9��gc��f��bL��^��im��,g���[4P_[�hK<GC��o,$�Q�*�Ci�t�SbgwU��T�G�?���%�/ԙ�I�������)��Z������^ mAX�z�P���2-�	j�ICs�f[=ɤ�&U?�����j�T�'@@mOU�!�
#��4��qIF]��/�O�D(���JkJ��2�	D�*������J݄��R�U*��8q)���}�K�3^"|4|���a�}�����U ��t�'�����;��CQː3m��$�#��w��Z�ZR���Q`֕O�+��)�����$^�_ꏓ����F��p�Ł=�<#�����,ƫ�h�D�R�ӣ��+l{R����):h3$䇤w�3�{�A�vKˍɘ�.��J��"\�]��x�r;� r���k�V�rR#����l�Q�XQ�g	Am��E��9l}�PߕY��z6ca#����i�!�:��]+~@����lx���O�<�9�	Nٴr��N#y�ɨ��dp�9��������OL4m��S����ff������<� �f$���c��E\6%���n@;���GfΉVc��>D���W�[�{-3Ndwm.�別��	�� ���;���Z�;�y�^>n���t����lƥa�+%����i>��^�t��u1y/���/>)�At�:~D�x�7��}�tI���g��I��%����5i�ݖ$�v����专�X�֕{����jn�ư�PD��yG*M�1�^���"|�`����bF7_M{k��n�b�,'؃>�d��L7F�'jJ�DZ���i����Ŝ�t�N8~�:�/N%�N�c��y�?�T�;�K��Û�l�tg�E�߫��{�<��U��[g}�o���
\)K�~� u@7��q.%��!��U��&#a��-@��b�O'ۑ�r�N�� �|����lq�l�ff3J� #�N]�<��h�ׯ-�ßr��y��f{�=��V~��:1�hu��THa�~2$�5/wOyi-���Z�Bi���!��� wBF�+���_ŕ '7�+M��2s��T߷�.�k��n>s;�dX��O1�5G.*���Ծq'�8Z�4��)k����7�N٣�y�p�K��F�!�=��n��H������9��F�a�3��"�Q��u�4���WܢX��o��LyEϭ�Y�ٻ�u�pju���}F�}�����9jWL���*���-$�*9��{���:�p�e���o���q-m��Ё��Tb����n[�I8F����޽��/P�h�"�'�_����#�	�m�.�G9@�nF��^��ч��h/�tsm�h��7�J��B*��4H�2?��t�.y��*K������?9?�b��,)��f����W��9C�P��eWuBC*����6�!��^C���S���lȉ:� �&_�� ��Ҟш��G���S�(|���O&!��0�J�@�ܞq�9��a7cBW$&]\�ќ��^(8�I2���9���;3z�4%T�}!��?&z1.����4F˒Q��t��T}���!��8+����^\�~�l��%U�LR��^3�5�����{��j�N7~4y���4����2=�:9<?���ymx�3W+�[}��{m�/�k]��6���;\d�DS��_�H������8�O �ͩ5���Ϥ^�"z�VVwʞ�«�f*�&:�]�r8|zJ2���rw������<}~0��Y9�<����q�y�����r?é.���w�<8v���He�n��цjq����y���	��6����ȝQY����_�L���D�W�-�e��Zض��&�ӏ�N���x5��*z4�-O�
c���9�%�S��E?��K�[g�bm�)K�VE˯���߈�j��rs���&�n]M�����	��$}>֟�Zlq��hP!rq�lk��/N�W��Q�0��E��oe�Ze�[%x��b�u��a~d�xRh��r��0��$)�����M��I�3����zp�R��vppZ��"��Sm�$R,c�ʾ
�}�s ��Ц(ҪN=\�
���@@`�Y� ���'�_�W��B�^��M�#��ވ~	��;����7�H��V�����ۏ�{fFq�K�
�0�0��V�"��(��������Y��"�]���`:�3unO2u�B�d����~Ond5#z�|atn4ș���Z��W��%1sC�_֌�Mdnz�jh운-c4G��:��AHC�ES=+�0�s0�mR�}TJݫ
?;�R�P�r�<^W��>[vY.^���i6��mz,]���ڟM�;��	��j��,ɘ$W7hF�N��=��_Km�\q����껅xx���cA�����
�8�O��ChZ6L�n�7\�(��.G;3&!��e�a"о$��0"1�C4����-d�MO�l,NB�&���\��+d:3�S��P��ۼ�7����|��a[�]:Y� ͒&���id*F���&�ćfN�Q��i��/�?H�s@��)���oI`:f�V���XD�}F}s\ɦI�P�v����<])�-z.*����,#;i�J�1o1���7�_G:�"�E��*h�9�zG�!p��=�W��B;��/����d�x��o�:q�Y�YE�:T�m�[��'$�՚�W���iPt���P�Y}�N�]�r
���$4�2d���2J�M��0*'"���h�P'1�-$a"0lc'>K�{�SK`��C`�껂�K���Lo���>��{��ҥ�|�h&I����������
��ŕa���u4�l��w/�/�GQ�����5�)"���1��/�9�?I�oxK�� Zً�U�
a��y�zZ��F�y���C<�2x�t�\����`"�_��6gP��w���:N	�s���� =H�6�F	�$6�6��
�f�[R#��}gy@�f5��ģk�G������k�J� �j�(�����")����3=t�n6���6�Q���lo��Z�T�����#1�D���b�:� c�q`��sl��tW�V03���aJ���?���l��DĨn6�p�mݺ�$C���p��ޖH� ���n�
rǴ��eN��L	<��c ����y3�m'�X�U��9�3_g#pE�m�Js�����۶z��1���ؠ,����h��}��Q�0��8�x�	�ڃ,�k�Ӂ9k\`̅�s����N�rO��r�$x���ƽ��V��6����#>�D�Z�B�о��8/���VW��33��;@2?�/�r�:\�s��U0�S}����9O��
�tEm�#=S�#��T�\��o%���"�a}�/�PA���[���ZF�F0-\��i7�qO%�����;/Ky������C�Y}��з�lA`��.�Uj�fx�W�%�
�@k	ql��Q�����%6b��6���M�h�86xő(�l�9H��u��-�"�ׁ[Oi�@�5�b�z�Q�f�T_<>߲��g�Z��6�
R�*IP������2�0��Z���k�m．���tb���E����ȑlm� �˚��֕j�-9%�0�W��uͯq����'BM�Q��k�h[/���w�)?�6&��h��˜<��t�{+�]/�N*�H�gr�Ts�^`OØ%
 z+c�}�{%�ϙo3H�=Ke��$2�ROS�ǝ�i��*�}�"�<S�RQKp����Ϛu.��kz�Q'�|���O\~vp�t&Ҋ���tT#�bsF�cz���A�-�d�`�ı;�L�!�n�g�|̗0@��(ͧS�ƅ���-:Cwm0���^݌_'�\�>�L�x��L�����7�>6b�w�=Ӟx�%��t���.R����M4�$]|lI�nrZmB@I��hn1:V� �|0,�^�Lu�5	\i�N�O�.���nT�
.�mY�I�G��i_� dN=��<�?d��3J��LR\��>(�h�.�v-���12mR�S��|4�a ��p�K�f�V�p�6���L_�}��w��L�[8�Eʴ	�=�B�(	U�Y@��;V�՗�4�rJ�� ��-�,<�$�0�dO�NG���"�ȳ�Y����� >�-���;�i������)-�݋y^��U�5	�vtQ�<}9EA������k�I�=O���?���̪V���k4(��=	�{!z쀍����{=>����^U(��1�ޯ�fV4��1B��i�W�(�>����3�|y�������_��k�͓-Gz��ZтFD�c��w�Ҝ�v�0��E���`&�[(w���h�a��*�ȼ��J��b?��QZU���[_tӀ�8��;���%~
��ӉLg��?�\�46�Qv�QrQXL�w��)$$��,I��HHdʞ4�`���J�����m~�`S��~QAm�𠻎�k6$q���d�}M	� RO1�*�n�F�Y��b�Qy����5�����?� O�<��N�fc�&S�5y��Y�^�'Y}Z��G�Ui�EM
���nv���B�J�=8��Ѭ�lA�S��x���)���xҐ�w�Q{�5��bX�f�á�Fr]N����T�h��k;$㈇��53Aj9�D	�0@1}&5¨Ww���oɨ7�=��0�C
�Uy����s�xs=��lz��Ky)�h�����st�f���賑��C;$��N� ?��YTZ��!Yb*OG7z��p9�$k*�VE.�������t��x�W�����@pI`�zV${>�U�ؽ�3�w_��.��\
�`��8z���q��.� ��gn�t�[��.�曎�*y�FЅRj{T3�r����nRRh����î�܆kB`)�ᛗ��/�r'G�<&�ݡg�;�*�<����!������j�c�����R�8�zX\�i�`�fFT�˝=7��;�7� �ѹ��	��{ g�#fht5[R_�7D��hٮ*�?���A%@�4U��/^������_��X5�&Sp�٢Q���6<�3��Gak�r�F�4��ye�YeK�8&��0���N���X,t�h����fȵ+�'CȦ����f��'��uh.D�Qu�����3���M�w4?���ɓ��k��y~x�t�w&V��T��P͉�C<s ()6�˥	�����'��vU�X�l��,�#����\d��o��k�Q*�������s�c�G���p�� �1����i.�ޝ5���y�)/�����3���Ez6n� ����
��	K'@^�ҧ*ܝۻ��˛�[T�|xn��D L��}�Y��X"/1;l�`�5]�E�
lns.�[:5�y ���ɥ�&ؖ�� t��e�C��Quk��ﰨ���b�y�L�5s���Qh'�S>U'F�x�LK��� AnV���>��4���-�!�H鷐��j��[!X��i��ގZ���M�>����� �<1&��wR|�9�9����ȏ�>� K☐�����D`�d��u$���j����02�����3�}���;;>p)/�{�]�Hb�l
�]%F�����Ize�8�}lvU���j������+�d����C�%i%�����@j2�F�L2�،����z��}�i���+�E�?��̎h���A]A��Ϸ�8e6,U��SwBe�X�B�O�M���ޢ�;l�h}�}���;�:��I@{�,{�Mu
c䉡���i2����C�41,j�$��n�7�Q���O��$���K9��a����L���i��)��P���Kf�-� �9e�f"L���1]��~���8<����P�&Ն=T��<���AԐ�lA$l@��J�~��S*[��;��J|��ȴ`��LN :$hC�r |������	��ϋ�p ��@YFdm["OPV~,������?H,BL���Q�����Z��	Im�tc��G&:�EAz�wG�^���<D��Y��$�r{���V�15�ؙH��n	c��� g>՜�4S(����0�P�N6R��Z���)D���WF�ڨ�?-z�@��g|E�ҁ,]2��Q?K����}��XH���>�j,�����j\̐O�J?H�lw�5@���&七g����c�}[H�+9:��o�=�2���^.2��ټ��͙�b�dh�dU=��*�	��#\�H�Rtn�h��?��Ι�s#��T,�1֎�	m¤B�o	_#j(Ƀ�Fthf�9���2s��7+-�@
J��UQ�Gc���U3�T��@�?'��nG�h���i�/M�ҏkQ�2qG�`�?���� ���tU���T��/}@��E�DӹKz�o����$"o��櫾愈���5��!�'��ܴ���]u���.�9/��~F�md,MƇ
��uB�}A/�R9%��Xx�P��|�T0hGn�{�S�ij�Mp��@隶�á?hK`�Q������Bm��jIss��3j_�Ƣ3���7��d
�L�ƿaUB�!�a�Ou�T��d�8��e���0�gW;��v��1��� ��^X<Q�^D-��G5��J������g�	W��B�"ѸP��yy=B���G�<#QHC��>L���
����������(ѝ�k�2����ȫ����CI1P�Cy���
ys��l����&IhL��kf�����l��hz*sҧ�iZi�B���Qu��Mc$����miZ��|��KŀZ&6��^�Mfu�;�ʫ������p��%ZY�-2p�F�3�Bj��d��D}j�G�U���E�	�UצgB�"$Tr�8�d�8��
��3ؔ��cXk�D���'��+{Z
6j�2F.z'a��N�"q:s$������e[�[�YqN�t������F������Ƙ��iM����c��х��эD-o	�x)�a��2���m0�b�B�*T��1@�5@����V�Rz�y�%!�e^H&$��7BN��9X��e -����G�a�؆6�U�2��:�,{t�#�W*ggT�v4V�'�F��Gw-��\Q;���Z���z�*{�AX�)(�A�gC<�����G}�qv��;\k{啽}�n��_�x9��=���/�|r�{�_2�i`g�O����1+�轭{CL�3��� Lyd:��/���y;��3U���H��d��V����C�D���|��O��x�Vh�6�X��[�Z�;.�8.��T����A��>��(�+�gH�͝h����4���p�$o}5�M��59��s�͓���P~�f������::	��?�FWIݾ��_Gt�1�yt���j� �~��G.s���RȻ�'b� �������h�-'�H<\ٶ���m��G�9�6���C�`�����^�n��*I�}�uAL���Vt'fW��%�f��@פ��Y��������X��N���%��6p"Fe��2�����;�_z�!4с-���P��5��b��V����z�4x��.��ŧ�U}����uq�짙�ӈm��<7k�F�MIe�����W.�x�ai�\:_E�:���m�-�[W��
�pÂ���"�ZȒ`��ޫ$������
�S�.8جzR��]Ƒ������£НVwWW�/=H��*8��ޛ��K�(����l�E���4��#v��x��p��:� �.ޛ=U�.t��fVSLt��>�M�Nl�N�������y���ޜ�#��[<"[���G�*����2Q�S��䦠�~�*��C���Yڮ�3ߐ����)�C�C���	,ȹ�s�qÆI��&r���=���)`�M懀x�Lc�z5���֡���u��N����W:*���T];]X��Q �6�C��ߜ�2Ll�R�lJXY�y�s�.?AoR����@���P�^?��t�p�V�)�9��E�9�d<s�>����f~����92,S���BE��/	��M��Q�jם[X��'��8�~��T%x;�����q���\�D�ձY��v�����֭���kC4��ߏ5i�������/��.-7��'�}!~�#ûy3��a�|�C>�D���h�`E�ϟ�*���4�v:��^��l�Ђ��HJ)�8o�����e�;ќ��(K�SCX�]$�{�)��,����e�r���o۸A����_s��s���ޫ�ղs�'���*-���l�82[��i�&�\�<8%v�؟zuv;��L�S>����[𐢌37?D]Ss"nK2�z.��G����>R��+�]�"آ���î�(����Ta�����ә�[���x�;�[H��%y��W$HqVVߢ�_X%��Z4��=���@;��h��Pb��Sd�讂[áOcj7븝;�bVba.��1e{�ڄ$Y]�B<��	�w'�IO�t�#_�LP�v��8h?�Q\Ht�qPJ�����V�@њ0�P�p��/��J�����S&H�G?Z��t�}:���9n<]�l�0��8|co%H:+��P�6�y��Œ�ƣ�4�.�hxC_��&�ڒVm1Y��}2;n���("��	���Hf��Ӈ��_�2$��C��P���2��1>f�CM��/�d��Q��I��r&e�&�Nu.q�E'�����������+E��z'?ĺ�����n�E�0͔��9���`�����GM`Z��B�Eb/-#�7�EP���kئ&7���ָP�xB�*�F������a{�q3�"���n'�(Ll���s�F�H�kÚ�JF�J��^�����*5do�:�H*bQ�O��S�S��:�R�v��F��K_o���REN�A��M��i�C��X 4��hH�"�8sF5qڬ�K�Mm�G}�+�`<����V9Z���D�')��zB��"赅�ɍ'���l{������Kv�A\Tǽ�^P�@�Nn�
"��F]kBS.wխl,���u��-�n��$.�̠�����������K���Q����L�����
^/��/&��~�FPM���o�OH��}��հ�Nr �k��XY�q����2�|:�'�>4a@�]#ՑW�z9;�BZF��y�B�	���$��K�J�,�~"�w�_�y}�2Q"r�h6g�:ɞs5����<ܑ�I �8�n��8ב�_b����Q���ה���xލ�,K;#�)�8|?�RR �F�������Ql>4��i	'��;4����1X�iDT{�m����"{���y�̘�te���(���ݾ�e�a����F�Iǐ� �'������C����H��n���Od:w�|ט�V�'�0L��l��_+��8a��q�E	L~�so����J�������2���cRQ)�X�5"�+�l�Z�[��.�vT��j{Lw@�>���dG}�Y8�;����Fm�HS����x��1,R�� i�-����1��pO`��?d�`�C��y̉�&��8?D�k)�-��g����1K�T�@(�|���(ڋA����5M"-aֲF]yy2Z�j�a?8��2B�d*}����h����2�VG�1�_Z`�OӲ��< ������G�s����e&`�b�e��nѼ������ ����j�A�fve���V�`�"�cНnn~��	jWT)�~�PXPO�kfÙ-�����5���c�ߓ�AFJ����o��4cz���i��
�����={����T�su�˽���&��l��C)J̓!��R�>��<��%/���_OY�F���'��{Í���͞�uq���r�$�y��ࣶUd��<��|��`��r��1�n�NH��a�_��!�I�b���o��z�
cK�_3�_?�z�W�%�p��a@Z�ԓ�!*y��Z�bK/p���Z���tn�@!�H��������C����Xءr��p��D�E�s/f>@���c��c��>&Og�*��C�Yr��K�������͙��9[,�����B9l���W0_^�`��U�[�h�?�kl�(���]�����!�����������h��p`:�Ze���IX�/A�&,'��ޞ��.� ������Kb��D��2ސ:��&��<1~����SB\z�'����dq��澖$�<K=�)E����k//F
y��8G�+�j�D�)7��`��-8cGG�n� lGϳ"E��]>�[���q��'CQ�?FY���`���ө/b?ά�}X���g(�Q�����U�
�<����ʚY�ߴ^~����hb_jONT㙞%]�=��j����O[@rqy��s��e�͏ 4<�
O.Z���&�j��!t_݆��*ͦ䄡�E�ط�r��c+�����/�Ql;"�`��H�zn��=ܩ~̐w1�a�혓���Q��J	땸��	�@+ڟ�Xt45I�{�����yQ$��Ku0�w�텪��֒�M�b�N�ؾ���<���{-�>*�
&*�2JU-�_T�$�����$܂�)4_�,����Hҽ��l�q�,O�O�Q�e�Rj*6��ڥx��N܄.?-,���S_`#2��r̕"���)�)��:$�^��݊nlð���A��Y�!(��]�N`�<ݗ!�ʖ0
e���=�eY��"~B2���7�f��ȩ��.W��"໏���%�č��7��+H_W��|�zj�D*��%��QJ�C-�=�@�p�Ki��?k�3�W�F��o�+|#�P �kcc�}�����r2�4�P:+'5F�$��MH��P��Ć|������CMU�NC�V( 8�ޗY���'��
 Pc�q�7�~�����
f�'��-%P<;���� L�g+��"�m�K�D����[5�⃨ZB�ϟ�� ��`v��;�0��;�],��x��;A�R-]�?|�����N��*���+-�x��y����� qD&f3���]�ٴ�W#��N�}ͼ���]%��2_پM3D���L1%��s��%ݽ��7�C��)�i	��6Dh8��G�h�r�\�2�jJ9
+��ހu��eM���0��Oo�l���>UX�gQ*���,�ݶ {JV��zR�B�E�j;��q�Mn�*�j�������k�g7�2�'��rd^r�|r�l�N����3�a�}�d.�W�?�9��eQ�ɟ9Rq5�jV�F%��F�!��n5���P{X�Kx�BU��&J�E�ˣ�
҂����1����L�:::� �\y4X�nΎX�L�po*���~�=nk�ŵ�C��C�/�"��ŀutq �����[p+���Iq���N��UN��|;w�j�']��v���IH!m�*�3�C������s<����� �$E"��pm��b�cJU��{I��y-�g��5k�cw�9�Z�5}���럺�<�t��[1��ß���{�!��|�t�12���%]�xGNw���D��r���T*c��%T]�> y.�,��\�O@$�e"���\��"%�r����5�kv�C��β����P���p�"��D���_'e��O��k���v8T���R�����8��� ��R]J�A0�.��J�͹ʚf����d/�C�#&��mAFU�v�����6�Cѥ�Ygt���L�q������\]�؉���*��TڞD�r�p����5�=|����IR�w�H#u��.0U���~�`(�G(��!nғ&���k�7�pN��������8ql�Ss����߯��|Ź�9�8Z�|N�����HBDSv��B�]��!��1�+8�`;F)���	��j�X"]�
`MX?ӥgd�w���M�K��E<�R���h�(t��QAN!Ax51�L}�l��3�+Ӌ���>yĲ�F�����/!��&�W�*�N��IktŇ*>�E�˝J�Zg��e��B�����2����8���e�1n{��)I�G�R���:��z^!�p{ = ���i�d)uRՊH>J�*[�C�o���}�$ќ�4�����r�Z�>��2��}D�~���$.���-�3�6��;j�`-��&4c$��g27m�ۺ]�N�);��O��ᆳ�;�"`ٔ�(̐�����5gB�V��VYQQw,H�LU�&���h��݂�d��fK�����-#�M?E(r��U��g؏s~�L�kX�Y��ȟ2K� �JcZ�4�@�W7��~"�mS���V꥘����%�$���ft/��w����f�2��{�a�  ��@�W6�ݥ�^��	&�W�����:V��\�2g7�k��c�[K���yV�����y%�w2%1��`�����i��$߻��L�e�X3X�:<ȣ��ܮ���j�X����E������;9���c�Gs�,�7a��AZ�
�.����̿;��1�d�D����N�\]����&]5�������
�2v�n����2�M+p����Y�E�� D��5��h�̠�Th<�r;U�e���SJ�YEkl~��5D�����/0��E�{���(�h1�ܐ�J���h��N������]�W�v��
b�,�=�I)�n�����[>��I�Xyn��G�_����WH����=�j������)����3�0�G��ʅ{��p�J-׶Np_nl$|�CV�RT9�1CB�u*�	[�;|�����֏��m�4ũey�p��a����h.:� �����ߴo��u�A��
�:5?��!�;���^��=��.����B)����:jj��Y�-uE�����E
u��ks�3l�H�-��9*��с�0N�RCX�3�0�Ȍ7�3�X|5�O��{H��{4����(Vm�({c�g�1�FI�%L�b�
9�H�ȣI<	���~d/U�{�����Rk���[k�UM�3�^ڟ4�u)�޵�AԿ�ϗ2���7j��_ȗػ�Z��/.�=��p����nm���S�&^h�8\�p {xy*���P��Thآ���dgщ�~4�xY�ˀ���;ɯ�%�����d�YiA{�Q<��۾=A��h~`�gƽE�G���-x����<�p=��o�&�'��14au���B]P�1H��O�����#�s�ƽHxr'�?�kqP=��	U�tkPʭ�	z�H�%��.:�5�rT6|�u�bkm��t/L�W�ˍ��t�	Ug�����Х�����0R!�;�?�Y��ܸ��9�)2h�:����B{��00Ե���	�������{��VT0���2����n�����LН(Xv�r�O�j:_�<6��7���:��Ŏ1o�&9z��D�����]a�ٿ�U4�gO@p���[W
�p��[P����ϙ�"�0�r��;���(>ӻ ,%?>��~�$Ѡh�^�8�8^2����*��\���I�|0x�D:S-����#�`Ln�ߥ"<H?��� `)�k��f�m�={5�uR/����0�ד��3�H
W��q�	�J�d/v��bm�mȂӦ�$�{�$�žy���]9���f߉;��YTC�Ԅn��$Å��-6�?���� _=%ՠ*1�b�,;��8�%&����	�pD��IG(�y�yϗ�D̘ �Z!!``Y�"_�VXOrn&������8����0�Ɗ9����%LY��SG�����a����1����H��ː�h�``e��&a=��rWaZ�����.:�/����3&<w��rSce��UI�e�`�?�h�g��a!�����hWhY�F�z�R�ts��q���S�2F���H	�[@muWRkq��v�u�
@v� ���༰eHtǖ��0���O,��!t@b��W���cU�'��Y��@��j��E���7�+���� �}Y!��6ջ��W̢���-jH�TJ~��_�.��
*�h1��h�g��tEV������PR���xܽ�%���(-`˄'_��L�L�!�܌͂���r�~f|�j�n׈�?9ڒu��3�@���1,Z�Cɏ
�-V$%���y����kü�p1���5�����y�M�O�l�?���l:�� �����i��XK�1p�oE&VBw�Ff}��� �\�����:��*,���~w?�߻.��{*7١��6l��|��`( ��sA�q�l�T/�HQ��O��r�f�N˷����~��^��%�ONG���=V� �gg;U �F���0�������W�%�PwGCAt�{7'Ow?n/ļ��=}�����ox������k@~��γ���vo����{Ff<�IV��ʩ���@6��G�&v�s���F���kl�9������Jk���ޙ��y����t{�n��1�=	/,�k�� �h�IG���[m@��|xp��5\K0%qC4n��k��L��ӗ�AX����e�f{�.)��>���/݇�N~��(���"��-$�,l�����Z3X����E��nK;V:���O	5g�yv�˝�$����̸;��a��g���bەJ�3U�������Mn�U�������<C���7*��ж�v]�ϿX��{�Xy`�ۗ�!#j~�D�r�0~S���q�QE=�(��O=��ղQ�|�A�W(�yg��Y��=;U=q�b���M�^�;G<�p0?�����*���m������cE�W��A�d�HqI����
�s�$��>G'zz}�Lz����"���c�
�0yɽ�܊�`j;*2�b��!�ƞ�`���=V ��f-Ïz3
h��C�]I�,��-�1�5����$�(2�Gm!ͩ�;�+��e�6ݜ��~)H�g�J���v��������D�q�Y87|Ć}�tK��f�ό� Ũ�{/&`�'��-�4h���T�����!��U�k��>�M�sl�3a�Gu���@^τ��Ȁ�"�ȎQ�ᖌbI��+/F�`�.�����u�Wk{Dk<6}]z��]���g�Zt�B��"�B�s�c;zLd��7_�6_K��*}�`��[����!Z7��&O�a	w��B�V�M�Sb+�ڴ,*)@�9-�g}���.�(ӳ�8f�0�/Q!���k��i>K��w�6�󚆿X�Z��i��c+�����/϶�=�8��X��,iK�+}�J���B��/��h/�S�]!�h6�H�ꡐS����+����g3t�i� i���F�ټ�}"o�pxU�[�3�?�d}s��]M�`:Skt�}�&���xP���� w��ާ��F�l��{�͚X_��X+_��#�=��|$�n���|����ͅb;*���/`b=�P��辍	|W�	:�Sl�]�)=0�]Z@�"����Ñ��|n�ڀ�4�/.*��T:1�{��8���ZL�P'(�7��Q�)���pYE�C����άe��������X�t��t~P%�P� v�Oʻ��|���%4.��2����*�
���#\x$�����<��Ϸ�U���J*��IFa��=X�q�r�b���I�{:�Ұ:��`nMo��~��B�N����h�@�7�F|�MN:����l=y�C4��dh��<��D��l���]Yzc�6
����'r/Eu� �`#q���A�����v2w�BM ����L?Vm��q��͡�� ��_��.EW�D�2����?:l;��/�v]_�{�4��%�ߩ3�:�1��l��P�t�,�+�B(�3-j�j�s�E�*���A]��x��A�
�N����s�[����%3���Q#m0�@��ᬚ`�_y��N\��M�~���J���F裂����؊,.�G$��T��%�҉[~1G O_%p_˴|��t�_�%�|�<F���K��q4����b%HTKcZ����l�$.K���jF��Q�f��ȓzN�d�y�^Y���V���fT��~�0h��ހq�b� Ӻ*�R+� C*�&��g�ݿ�PƁ�sW�~%'qy�ҝ�"ܟVq��F]��.u�Z-j�$�s�W���J���\x�H�|�I��l׀d�i�r;=hds��z�ɟ��Y��'�8D1h?y�Bs�u�s�Vi��N�nJ�e�K~�B�JS����~ւZXs�R[Ṉ��I6��'�c�Ì7�QQ�v�bǠ&��~�~�����V�{��g�\�G����Q����l�5&�V�Q�
r�>S")�lɝLj��U�x���ͲV���*o�
�$���Ш�\�� �Vi��@�o�+������/�D)�Ѵпm0��@��֞s����b��X�fR��%��e���J��W:�b�|hز��w/�.�BP}:��[2=9-�B��P{j���i{��@��V��(�x ��Z�����`������H����ܔ�U��	��>?<T�N�Z�"������71Ԕ	n⟏ˣɇ"\���P��>(����h-��Ľ��������*��B�+���xH���.ʮ~�^�b�R�٘��$B���U��
r���*��c܇Ͼ�$�6B�a���w��z�O��u����&+XD��~R� �r"��hl{��U4���z'�g���u�l�/8R��H{�iO7Z��_�A��1�OT�J�6�G�,�#��TDɎ��+���Nsj�U�v3h=�k*&���.�Aj���r��lIZ!�����%�Gn(�X����j�]	��~��a��R�9��nX���i�Q�|�Y����p��� %��K�������f$yS��Ʀ��dz]C{�@�(�,)2��ր�W��c�Я��?����!��(˚zU�C w��S����w`���0�P�g�e� ���� 44cr�m^�z���Ώ�z&��_�
<�);����[���똆C�x��������1���P�|�d�Gm7��f$?k�*?�?��6s�a�Б2�P�S�ӒT�WoW����(^Ƞ�i��������F0��e�v�qS�ټwA�b����� ��̔�2��ׇ���?�ԳY�@|Gg+ ��-w~o�
��(&���&�xg@�e��9FkH��͙���VtѼ~8�\C��".}�Xe��'�vt�C��zN	�C ���o��g�*��٭ؔ�ig>�;�H�� �>-}�i��x��f�EzLq)L�w�[ @ShR��COD/8�/����?%f�����m��V��k
 ���0�a��ma<e�RΖ���Y�P�ȉ�2��C��5��׎�� f2f; `)ቇYޜQ/��M�6�V���(�bM%c+���XB8Z�S@97��k��Z'0��^�"�,��<Jӑ�{|����e���*L؊F�,�Añ��<ټ���įX<�/�����`�9�J���<��P�/%)1;���_VG�&���s���d�aԐ�rH�)U"�n�tK��,R_�7�b򈬍��"�ڞ`
ǿ���:��0�\\/Ǿ�!��PX��h�~���˻F���(&W��V̮N���qa��vքo?�������0S�ZE���b�:B�����q��k� �ǭ[U\����m��`�.BbY�v��֊�8y2���i�/�ː_Nr9H(-�x��r��'-Z\~6Qoؽ�h��,���(:����"5��eR����$��en��Ar&a�̓��-'�]֧�n%*6�%�a�!�H-���G�	"��L�I'Kj���9��m��D�5��:�\P�}w~�<�K��h�N�4j�IA*d�~cy��0�����	c�M0�2l7�O�U�����]˂������4x'`�� �-�H�u�O��V3�+��Ɲ�DJ�y�I{,�n��`	���Hi��pD�f𬬩��s [)�E�~_(X�s�]��@�Obկ~v�(�K�U]2�9W�����V�8�6%�O�!]D1���Й�m�Bs�'L�+"!۬���h���6ע �>E�F�����֌��Q=>#ӵ'��)]�`M�J5-����m;ƽbŠC�o��:UލC��� ��U��+`���쏡��D"$9�l�%�c��Ւp���}G��g�J��Rh�T7�K��)5~�M��r��o7�5���K�_F+�#�шq�^<W���&��㸂үm��a���v���;�EKP�����h jL�ts�`�U�] %0羯}��/urfg�?����+(܀��;�\Xkç>�vfi�9�0�l|h7P�,a�V���]IP���kypl�̵h2B�6Zɟ��5��yyI��#����j~����ќЪ@�J�l*�U�O�#L�����F�J���M$
��c�����[ku�����d�e����TŊ�
Ǹ�o|����(y���G��N8���{a��b���*���vbG0.4��5ϽW��lt�u�M�n�
o���U'� ��1�랑ۑ�]k��(��zNC�$x ���7��wn��Î�M�6�R������E���ބ���J�{ �]Y���#Ҥ�F��vJ��E2��94��eU�9U?���t:Y��:��������D�
��#BSTvu.��Go�4�cs
}���kbv�R�X��5��pA���ᣴߍr/�0dG����Kc1M�5��@�T���:�1֘+��M���!Hv���Xoyx,S�!._/�ms�,p��Wc�! ~M*��"���)�Y���d<sǑ���ޖ?J��Q�~�^tgD:�2x`q]O~��9:߬ź���'��Y�fyCT�&?<���
Z��o yɪ����נϮE�0
H &g�/��Z��SC��ld/څlM̓�1	��pD���kMݓ��D*�G3N��ױlE �Q�Ap⑹���O5��$P"�a��&�ōL�;��'��7��UAQ�C���d!�=�0��R'�b����*�G�ԁ��*?r"��i���ۡx�ϥ��� �X�C+��슴b�Nt�s���c��+W�v^��g�)��R���E�-�j4���Q��p��{Z�k� !�lC�A�Bu��:�P�ޛ�*�A���ٷ�@®А@�P�7�>8a��aUf�EO.�؟�L�8>���Zx;چ��f���2��ڵ�N���酏*\=��j��[��^�����IR�Ƽ��0���Z�� ����6n2����n 3�[��{�K�3�:�冀�����ҹ��+_{�'���hU�ZC���D�ݒ��;m�P0���?歨�m��f�$-ЇyG^2�L�DVS�i��ҟ��Q��4���mnH�&q+� +ܕ��7����:?{�aE�i�̌��}CB��Ĝd���c��g�+�-M�zk�}��R#����J�u�_���.��o�V�����3�Խ�+H�Zf�/���Ј���nJ�{Gf|l�4���򕴗�k�,�lݦe��������� �5��A��% ڍD���p�>%�/��L ��T;|0sW~x>��ü)�z�]`�kM��[�a��\U�ͳ0�D�?��^d�һv����T�9𕱱.�-m<��v�t��)�Y��7� +W3�h]��]��cl��C�ֹѷ��@��\p4Ibf�sC���ux^�ƕ4Ug��h�n�Q,Y�����iޚ;�
���R���d�*�y����vX�+Y��>J�(��e��ǔ��S�N��h�8C?]k|�����(?���UTMHv?�5�c����� G
�c��¥��$����ѭ���Z/�Kﳏ� �Kr��C�,Ggo���� �[D�f���)���"��͹.��c8:��Ʉj�e�EQ��.��ȞU������[9Q���K%��$�C˛N7��K��C���a����	�V-��T�4S!�MA�~�}��_�D�/ȟ.x�K"���~���]�����(e��+�a���Q\�������Wf&?�����[J-(��
�nntHN��eϛ��k�Q�7���wt�����C�ق��ˉs�#�1j�s�� �H���T�/؀+�D���q�4��z~��:�Q��^ ȃq�u��M��1Nq�P$Hq�$�O�j�����By��*?l����<KRB8 )�������TO�1����3�T��q��m��2�R�]�xz��d�w,���L�FÌ��A��3d�F��ܲN�⎿��Z��tnwc >:�G������i��|��n�j��à�&Fh#_4��]���=aQ�o2��I���ɝ�(�W��AB]]���+Cz�H�E��3��4��q�l���s⁡|��Z�'���e4�����ԡ$��P݃.V���T^�<��[r�|'{�j�Ǒn}�9�v�b
�
�v�`K�Hz�C������L#�
[��]�qS7��o�Ћ����)��~V�r��2�+�[m�y�%�ײ ���o�X�(�mݗ���h`/"FK�Tq�|���x�\
T�7A�֡>N�f�<��jޔ�?�`
�"Z�9irݫݶ�8�N� ��9CL����8f����'Jg�q�̣\���������yYN�1�K�uN��S�a�8fE[5
L����SM)�=�k	t�`Q�wBAs!Zt��E��Pg.l�̠Mp���Dg8sગwV�b�������+LH�<G/2�¢�חר�7�3
����dh0rusF��(uAo��ْ7�%h�Rv�"�^s�d�x��$d�0IǮ��ܨ/�ʀb:w�@8�����I�I���^T�r*�չ��b��.��|�H���b�
���am��"7����ER�\
�D�Zd�j	����:�}
;c��&�K,�%�4�x60���b��#x2�"�)���y�[�."��߂Xs�n�φ/%����Y��1����L��.i��A��;?_�Rff�%�#����z��dY+���R5�QBY\�����z���]�,j���}�P�N��5ىڋN���o�h���G�̵g1/��>� zw`�8nfJ$�s�S^w9��C
A�=��}?貊��P�����^}=77ӵU`����꽪[�����$?�p�
H�����d�>�FO�.������Bk5��Nx?���TB�}��|T7Q�3ڭ�]v�xS+�ԏS-��螭�u��L�+�����2J���9s��9ؒl�B��O�
��\4��-S�xi���~}p��Zsk��~��>h1rf�ʺ���V�:GǚG���-߃��W<�T,X���G!w���Y+fm�������&w�4���)B	�]?��A��v��M���Cf�����E1C�t：�w��r���H�g��b_�**�8�	]���<�n����XW~���=��K�M���W�ˊ,D�)v�����Z�\r8�7��V����@m�-����'���r�����`g�k^��>�D���
����2�֕��܂�<X+�ehu�~�F�v֊0
2:�s��F��KU�U�b.q%��-_m���i��坺��բ2�fq�`z��zi���!���D�i��D���m�v�Ì���h�y0� ����v�۽酊�
�QC�I(i���K�zs��Q�YĊ.����z$�\o^�<kZ�~ Z��`V>Cά�/&t�1�����G��V����X4"�U
��b�Й�X�W����@��
�AʠH��}q��o��t���:4!П��d=�Qǰ����͸�N�P��1�lƕ�)d��K��6�ӆ9��GU5�փc���F���OC$>��]E��J��~�䓏�m���[7����q����RA��\'+ñ�8�.כ�[[�,������S5�#t��*�9�`/b�0�)�����~�=�R�Bn/[�{�ΧH��'*j����T�c��ԡ�s~ϐr��� 8� ��r*�*^&�%j�F�D����E�g�kܛ�K�E�����ӡTh����4SӼ�M2&�wf�p��T����K�<�����S�U*���3ee\�]/\�*X}z�@�]&��5裁�Q��ǟ-����U�Ykwx(�Ç���pRʗ�~�
��������Z!V�_����yE��犵\���C�b::S�O�H-Ś딂e��א�t2oa�^�{��K&�����"̫�`�T|��PxT���V�b�����(��]�1:>{��
�Ag�����7�<��������J�}��_� �O>���L>b�	a���{*��B����W�?��ZX���%ށ�5r�%[��Z�������m�A���W�]�@/_��V_D-��EozÆ~jU|��r�`�K�~�M?�]R�$o�,s2F8���v�i��&3;��Nz��I�L� ��7�mn��cORX_��;��s2�m�i���__7��R���E�+8�7�5}M==)Rz'�c��{]�@�q�i�H@�����Z��QSuX�)����v	�=c��M;�A�#m�*��\|0� ���.�������]�Ɇ:����t�s�+��N�i�l���>ˇl5h8z����R�m�)>ӎ!��=���`���n��Z���V{UՖ�BE�����݂d�R�Gv��ީ���Ł��a�G�6W��`�>�_r��?���.�=Ɋ�N��󩵄Q0���������̃s� �Ǐ�=y\�"�w����ED�Pf�^˅���D��DDB<l1>��,{e�E�g@���c�dH��f���*�l��'�)��O7�3�Blj�`��/�s?KA��JV�<X�̥�����+�^*��T����z�C�_(�{���f��������E]w�����8xf�����\H.ś���>؛CG���S�;�ݬ���R$Z�)���R�E�Ǥ[G.H@68�_GI���!Ǳ�b�}���3���˳ǠQ	�@d�@-�H�@2�N��Qm^�g�8t���
��}˸:����b|�>m#Ϳ��{n��1�Vg0>�	�{�����_��e��:W���ua���&2!7�(Z�		@z�Q|�;���Y�~�ZBy�2�d�"���o�����\��^���y&�ݖ^�i��d�6� �0��s��}7�JI6����!"�PL6u�W�W��/�sn��������d�JJ�O�	��`���R*�k@�H��<tx "���ucp�C[��:��� ��1�f\�+|����'7M�c�x�`��z9H�,�X�\��+�	�I��o�\���,o��K��d�΅�K��0yyt����}����J�Ѭۼ4���"�J��c{�>�ƴġޠ�����������Kځ�c�ڱ��U��#{x
8�ˋ����J����a�1,��Sؚ]AH*N����q���($�Z	��e9�nȢ5i�ʋk��?�e���GV}����Vt*��$��.J{�0H��&��W��L��M-h'�l�^5�P�R��
���-w�/�/�U�ۼ��] �C�#��>�|>�Ԍ4�0[i�r�W#GzV@����{��A,�a儰�DrȄ�rY��_H/3���Pd�N��1�q��v�oP�cz3�a#�o��mW��� /� {t2�����$��-���{?��gҴD��DQ����:<�i�C���X��B��97��f�@��/h~;N��FYuK� Z��jSY��I�@�pG���	�L`���J�]�={�^��!9��?�����Pt�@�DT�Ĥ:�c?��8�6ÊKs�k&�X��ʑ�PJVZ8E�݉a��ٝ��M6,�I	�am��8�BI$=[;����5�� <Z��R�����.f����V���� ���5t~���=V���]hPu?1�PF����V�HU�x#�'cB��C �B�*vT�rs%&�*�\p8��~�������i*�V��i�87ʡ�؜��q����Q��-����}i�/�;[����-&rd
��W3y�"y��(�E��]n9����H��o��F��@���B��S9�����X^�� �?��lf�R�ʜ�PC{�s�呻2��O�ڸ�?f��z��g	��y�M���K6�Դ���ز��K��wP�KgZ�:%��|Y��+�G�?0�@��a6�
%�gͫ��qca�L�$�@m��T)>ĳ�"W�)�A�B7��%�_�.������wFw�9aT'qzt���4��[`!D�xZ,�R��,�i~)$�I߄`Ʊ�t֌�WCP �X���l��s��`'�~�?�^������8
��)�
xM�<��^�_X�zKWg�|1�al�p�)?e4�Y
p!qmؾ�J��1�酠o��s�W��,u��b��>��8�o*�*�P=K��6���!��0(Ǭ4���ZQ���tj����qd�k�b��@f���z���nƄ0�ꈬ��R%$n	�����l���`���{���ͱ�e�:�L:�3B_-�gN6-+��>�.;2_�`L��͸/�U������ew��8�#��h7�`\�]J��������c6������9�����T,�~�׆�@�k,%.J¸���'�n�n�^N@ɢ�vz-�E��BT�ij%dK����&��" ��$Q��k>*�	��kT�$gj�b`>��/��'�%�6��s��-���3E��?�=�p��=̞s��.�U}*k��}5�=³������5/�.��󿆾�H�Gc�`2�{%4��G�ǳ5�F�2�W��f})#�+�f<]D��j��N�>��^vp�Qqr�[M��S�j|�+8LWe��Fm[����g�b>{���v��ƶ��	:�)�HL:��ke-�R�i��Q-.��%&���J�N�t2e�`j0C鑟�!yHC�z�Pf�d��譊'RY���
Bgw��3Z�!>xQT����a���r���D�	���s�����r���\�:�H(��sL	~D.~����&`ve��&仰s�C�t����C��f&��~!�ɟ�Წ��Mܐ�6�{e���L�vw�Q�?�49'��G�DL�&;ܼc�б��p�cٌ����(
�!�ЃD�y�*,O�/a�	$��Ii�޽��!~Y�S����JF�j6۵v�{�*���2<"(����&W�ii.7�&"����	B��5��k�מ-�l]X:+l�ۓ�˘GQ��I���|t�J��8�۫A�4�����?'ï�y}Bh�Z� T��oV�-�QO�#�X��1X��ZR	�\l�y��2�����j�T��[�iJ�&��%�|�ͧ��U� �q?N*��_8��z���������y,�0��q����y�y��r;_%��'�;����UY�\g�L�O!DX򉏒���A1�J��[��q��P�N~���1ײ1���ˢ(����L��t��:g��1�H�S�9�e��lQ��_���/������kk�L�t�� �	.���9> �~C+|�D:�Ϯjm�:��6/��&���0��S���	~
��x�G�&��P�M�����Lo��eu��Q)
>�A
��e�<�GE�"�����M�g�茎�Uo�7�_W�~������9��w����Mj���$���%��<ϐ��t{��D�`c���S��8+>9{+2�*��D�
��
_��;���v���W��A`ԗ�g��ج<��&�ů�L��TRk���dI�Te �|�C�z<j�{;��&'���Kh1V�, �"[�`ηM���+���j���d�s\��� >ӯD�ޛ���V������p-�i���p�0̸�P\%$J獓���'Q*�e����:!q��7�������yz�֘qV5��;���������-J��,����_���\�Tn�s䂴���<�pzRLE#��e��O�D���<�0 LՍ�B5�i�N���V��쑐8}{_Ȍ>-�`H4�x�
�6��[��ŋ?ߎ�q^RTޫ��&��6_/��9`����8�&�l�-h"6�B����Z�Y�d��rYٙ<�!����Szj��x)��Ku.�5Qg��WY�n�V[������Zؑ�v���1`���-z�ƻ\+�
�ه�'_����G�@*P�|;.]�7���	�Ihxȣ�&�y��~�7�������C���yZNK0=zԐ��t\Q�B9��٠��uw O��ag|rt�E�� k��Xn��҅�ﯨ�oԑgF��%���g���	�O�JL�5��"�dg���ӦTK���⠛�p�E&���+�����2��w��6TQ0c|�V��J��z���Hm6��h�H��啍����ҽ��	��ٵ��w�h�n�p�cn�>�.H=RL�[.$/k�$k��kaY��� 4���j9e�N������Gqh\tF��)`pb썙$x��v@l3�
���Y˴�~��)1e��3��K�)����P���&C��~��!�eC��kNg�~�ܣ�l#�C�U�m����M���W����� 4ORl;ON�B�*��
��r�=X Va��u�������8��KT��	�7���fj�e퐊8���Vvf�On���{�s5
����*pf��E�Z�C�r!x�+��OQ�`��V�˲��`{p ���Z����P�`��%���o:\���I��]�v�����[}(�sߕy��~�74;<I�S��Q)�N�w��� �C�RB:m��DÞ����T�x��`��v5�"|*cGư�0�LYkXZJi�Ud����%�n��Yx�n|�9kcpN	�4y�S{4��-������F�}�L������X��GDb\I��Pܿѱ�n�����7�N����"w�}�����N8�H�8��5蒰1�������q$�^�6\���"��E1�������w��1E�����6�L�[
�;|�D�s�]7�~<G���k�=k@hf�ãI�����L���aS9����A��ǃn�b�\�7�ԅC�/�Pj�?���G��@���o*�[1�cIB'7�J����7�8*�p�Ue� .D���[���ܬ�u�&/��lZ5��E��ټh��0ŰY�ɢA��h@�{~�- v���Q�%�Ƌ��;+�g_h��m�3qx����8G���������g���vل;����]{��D
^���Q�� �H�C���O������t"�*
��6F�"1z90���:wZ����.�t������%N��5 ��� $��G�?�*}����z���&+'�R�s������"J.�5�Ĭ�;F#�2sk���W$x'��6��[�ۧ����@]���^��XK��^U�ñ8��t ����
5|��<{6X���Bi�~9�[;�VF�B9�GB�6/g����8h���T�2����'Ғ��2f$���;�{��"����S�0У#q�Yq�}���քW�h��<�O�����e]�)�᪳�DS+���y>���eGt`�>Ekv��
|P�ޙdu(�4��'�>���I�=y����=^�/��.��ATk=�-�}2���Z*8�.6k�ٽ��~?n;�s7mW��˯lHB�+ �3��Y@$���ǎQ2����J?)ԧWfw���"�4F%�m=tk(:<��>�S��nY���� ��-7m��\�I�$�󞁘�=�t�t4KK���{�Ú��7Lj�|�e�Z8���b�襻�ʹ8��QI��Ar{�����1�������
�Ĥ�/m5b�s��J!Z�x�3�"��]�h�$�7��qE�1�lm(�P(̑uW�`3fJ�V�L�r�Ε���=Q\/�ʬ��B\�<�Ѿ&?	5�)�CO�`)R����������ǈY$�T�n<<�O���}��znL؆Ä�+Tr��j0γ+i��j}�S{�m4�̶̤;� PeL-|�i�	��Lu֢1�J׈䁶l���@��!���uҷ��nM� (�dj��e�S�>�#��R�~���h3+����W�@}�qc{���Ǽ�k��!W>!�y��/հ����T���${+�}���s	�	����8s��6�j�>�g�z�#��c��4��-�zb��+j���y�#mUx��
��r�T9�7Y/������˘�G�]x�ςէ�d�h~.B�2i�����k�麨���V��z�,U^f=��J��xߋ�\�F�b�!\?����8Ǜ>́�O�5e-�R��;'����w���J��	��ǴL��Y+=�weJ���\�\�ւ3K��@;����.�ξv�=[���ث�NdS�IW�PY(���pO��i�<�������frˊ��[Ŧ�������Y����^���ݛ�>��t��k!��<o6�5|*���F&���/����A`@ hC��g�W䤝��\��ce��	�b`�22����\?� \�Ԍ�b����4���?�q�QI�K���[��p��l#�?�2f�m.;�P�
���"���b�%@��Q�����G�L�[�B�0�>������χ�6�t�WlC��pp.�^PС�$����QoH��b��jv��7T�O0tF"2� T��,�����wD���z��������>^�jՓ̏Li~7��I�"R�H��\�*�S�}n��'�C6'XoF)�Ë5��!g��$�Usk �N=T�Lz�8�,�r�D�߀�L��{��� bE�V%�����G�S��Z��7V֜��XxY���W
z�ҳ��!<JX����|ݪ���Ҁ4B6�Z1J-��h���c���Eؖ���}[:���)L���8��[{�W--���\�:@������~�vtќ�f6�x�p�Zfi ��~�/������� �
aLLaUb�83\��1i5l|������+2�:	���B$(��G��2�%���n��ScnX/��BP�_���$�I(�h��D90w���RG�p7�Ĝ8iQ��L��*�����q2�l�o�^��=�'B�*0�S���tZ#��b�^���`Ƚe��A��G,��0L�0�P��?���zy�ץd*'��[J�#�hEBf�	7�T����$�|��0X�Y��F2�i�w�� KO��ƪ�l�3s
7�!����Ze���5������̸\ka�" cWe�#hS)�~��N��hR�g��'���� �,���Iِ����Y�C�v�z�VӖ���=�����9Z�o���Gd�P���k9nل��G���"s��wrϝ�S�_C���'��w�a@^v��*f�(嚼k$J�1\721oD�4����~�lgh���d���o��l�T=r�E�XW�� !���>��Ot���wYm	����s3rZ��C�c�C��P�
��3Lz)�>C��:���U$2(�+����"��� �A����\Hh5��	C�*���]��T�� �u�� t�3f�"�o�/E�: ���A	���������)��{�Gս6��2mťlQ; �{g^	Y�lD�yl~+�_p��-��1���o�O~���#�T��^�u+�]lAI���uFI4c"��ZS�_��@)vT�S_l��b��!�K�훜4.�іwA�m�"b�KL;�e1z�~�/x����N���Z8�o���Su��6e�^뚅��:b7�~�͓��34����!��'�\��}Q����$ҶJ�k�nj��j��j�yA��m��ĉl~/$���uW�B
ᾍ�n��x_x1W]<ξ���I����`? �^��Z�{-.���ץ��D�Pd�*xҲ�9^�� �����L����W�WI��K��� R^��M�5��UȻ�?ZHknƸ8"o���f��ĳ���h�̬Xr�(���,vl$=�Iih�����?A���9΄I�� ��c��j@�.�����w����G3�tj�7�"�k5ȡ$�T]u��l�����1W��l�qZ`cdn����U�u�!�� �=FXP�A7��*����M(s�pK����~�uz������	��~�ӡ�R<��g���-�BC��'��9 ���]�h��<a���$l<����E���1_��A:z"��2�[���-�+��l�3�T5ab�v�ږ���Ŭ����E}��R��7JH���bld�r/��M�A�+���̔)�48hlS�I�kC��{��R����Er@�"�1˷P1sѢ2g�_�1��wq���ߠ n���kql�ыؽ-�A9Nz��1I�[X��~N�� 'ɟ��[�q�Ŵ5�U�C��gM�xV�i�\�hUډ���Ϣ{&D!��r�c[�!u�%^ў�)�0��������6�t����k�����F8��~i�'�Gsv��PaZƣ�3����+�����Xqh6�e���K�
�߆���J�z���0��0w�{d ��/z'���x�͞��,�WЮ�[�yn����j.���i�%0,:�W�7��*R��� 1�/:��ڬo��rH��8H?N�SP8�Y�S�r��U�������`�?mk%.�/���~{�!f���}3�8���H��,ƔS֧ �:���g�=/2��ۯbJ��v�;7�j)5���3B��8p�di�YѮFO�H�* 0�������[�Q��QH�A7*U�����}|R�
i�����}z&�y7��}�hN���\��8!-��.i/��qL������6�A���W������;���Q=8Y�C�pdm�T���ر�J�?��ra�(\��l�sny' fҁuˠ�,o�_Qo䆴 �r,�	eD��lK��^ͤS1��ʣ.�����+~��e(�Md��u}=4ͼ5�J/�{G��3t J,�	��c�t+��XԉPźc�6��Zn��W��3���Q��Z�53o�O�鱈 �gv{q?E'㘖�!h���f\<�"m�|m����(�����U�d�=�"�$x� �!�?r�y4��@@��b��Ty��O�t�Ko������T8��]G,A-1GP@p�ӣ��܋��G�+�S`%_a���d�v>Y���J��t�(�DZD����g�l�߉��'#��*8W?�������Q���ĳH�o*EF֢a	D{�Y�vcg) H�ĒB���V�ǫ텽�?�;~�9��6�x�<*zb(���&q�s��ɯ��s�="~b�E"���p���J�V���#*T-�>zd~T���#�}�������k�2���pE@F�\ј�̃{'�*w�9ǻ�X���|ȵ�Gي�x�P���{m�p�N�s{M\f@0��0ס����T!��2��t�K��Y�n�W�Nǈ�Q�J;����ᘑj22�p��=`�7K�)�`�~�y���Xp��P��5��_LC]<`�\z��[+�;����<_����7�N�Zῂ)M��H��(��F�`���;J�E�?.��9o�r-�������IW} -i��j� B��1�-w�2���C�vV�ܡa�q�/5�q����š�I��n��*+(/�r�d���WQ�(]�^�C8)����k�ށ^u<#��0��僥����i%�8����"{$�p�3�/i]��ljӔ@��M�>��#��4u]���vXf��E��蔻d��v���[TV�@��#��붆B�
2 &r�
�h������Ÿ�)ya3����lC0�s(i���wX���Z�	Z��������M͕��%�%+�[�B`{%�)|�F��t5Pa��Q3��2^��; �c�jB@��3����/,:�>�����_w,�������m"�p�}�,��ᤗ��WXoe��������h����?m����D�HAL�����lSw�F7��ʒ�w�e�M���O�V/������ה"�d'��&���Rp/Q��2��/�����e�r�i���)���o��v�b��fG���N�)пn�����e4����7�wꗰ��������׉[��}�Ql=���=8��e�T�AZ���.W����|�*�g/�M�=����N�_��5���&��U~�7ި"���s�+RH�b�$B�g�t�7}��!�$۞z�k�Glcd<k������h�U���2�O��'Jv�?��t��G���ȟ�+.�Uټ�|�0�^���$������R�d{��fn�[��ml/̌�/�tt�0�����[���eC+����M�����:`!Z�"-����p����F^o�p$�⠅����դ���`v'%-�L��e�1G�y�^	�����ڮ������(�M�)�E��(Z��o/�DE`q�#��^+��\�1���3�����Ř
�J�r�k\$��$�L��{?�j�f��|�j�����dfpq�}ϖ?V}��w.���OG���1,8#���CE+�,�ȱ�ZՎL�y�����7���>B�Q��Tj�*��}�������
��X�,|XQFR�X��o�`�D�E��Z<���1����:�`g(%|�QY�&
c���%i8uұ�-�N�D�B6�~r^���F��i3k{^6;�:p�LŰ@{8��w�"k�C��Οr�<;@37��M|a���z�D�6��q�I�f��q�2��[��[Q=]9���س&�}���.QY�i+/�t�x�l�J|{�_Q���ۍ�_�1s�y���~���^���*.���M0Z_ZY'�V����FGF2�� ��w�:a��QKi&���{~؎���=��\0��o
9�:�|b�G1�{����MQ���N��8�wJ�r \�%޵Yv$f��yku� �n��̺� ����y.����/ٔ|H_ ��4��9�:hY{��z���>��4Qx��顽W�����YnJ��h�CNY�};���D�_��R��\ݢ�h��~��0��ހLO�� <�ꀧu�r
��
�a.󞍬����e6^jU�)��2Q�@'$(��/:�]�\���cc�!�W?U��-���~�c3�+=vڮ�j�����!��<�$��pF��"H*o�����ǲ�k�	���щq}Yi�**R���ϫ��������71�d��b��b��.�E|=��`�!#��>~��k1�D�p���>�q��E�D�V'nv��q��F��� '8O��	.^D8ǯ����\~��j���&u�2R48H�9��UN_��?��4��]��AS��U��}G�7�F���Yq\��p��"S������Ӓ�<k�Φ�*�Z�;�fN���#X�F��ʘ�c�I�z`��[Pr>f��}Ev���ul��i1X�m�(?bv�G �H/+Ԋp׭=�G�������G#p�I'�h3_�w"���^��5�M8a�S����ʓ�F4�n�C�i
�����{Z��Ģ7̔~�}� �H~o���9�G\x�A�Ԉ��0���"��Ez׿�bp<��	WJ,����N�o�fDo�b1]lj��y��B]J����^��=i�U�����!;�媿6�KZ]�n��65zʵ��]�$�;�?�=��=��6E�H�d��1p��z`̀�~e��=*�S��,�A�<䤫��W�'PΟ����b����T~��.���� �G(�Ѕ�k����v�K5�i�w�{�lrx{΁uO,�=��DJ�p5�ݫ3˩�:/Wm��I��*�&����I��SB=_6{ ���CH������6�5(\<f�yh�DPC|���~ؘ�o��q�@Ռ{�����Z	��V�mf;�v;�����M�+9D�~�v� ��r,�u��Ej�=�GuX�����N�f���8>�VAluY�/��j\8�O< �g~qU�m�bp�V[֐��������,��[L>J�{+r��wBa���D�]�$�����c�=yV��6��~��`[�$���07��M�6�w	���A�>U.�h���^�3}/�P��6b�Λ��v���\�,�A�x<l>�����j8+{�YLwh|���F)-'�i��ٲ�7�j!���Y��b����m�&+�10�M8�Z�8&ݟn+�����||E*Z�9�$����$Ҫ0)���X(��7���ժT#����.���N&BBء"������Jk}0||�-�<1��f_Cu����*3��wb��� ���F�Qh5�)�bM$,}H���Z˪�����(P}�~Q&ͦ��Vc����9��*��b;��ЭG�X��ٷ3+����K�8k|[f�QK���?��]8�����	Oe�9����%�1��c�=�A�����Ncñ���4�����S~���'��	��i_�r:{w�~�!Pp�M+������e��p�(p:n�<�+�����j-r+I���r���2����e/k����o'��Ż�tXzZ��ʐ�f��1;��ɳf���Q�bUylu*+�+����m_����+��oB��u��P�� �n���".!ۗW{d<U��$0|�G�7� @�Hb���C�&�����y���[>yXO9r*>��!�+��=�y��(�
$��UjLT�����ԟ���zA��X=���$A�f������TJ�V
5��=�������ra�d��Fi�3�K�q��͗����/�ֲr��aɣ"lp��t� ��Q�<�����3%���S(P���OA���B�8�N�ݛ�����i��J9��p	�U�>0��M��ۤrEA�y��<�����0��DlA��AG��Lw��5�hV� �����mq}č#&K���|�)I� z=bg\#kO�gĻ{����0��H��׬
w�0���ߔqL���`�9����h���фE�lט�E{D���)�v^��S�Z!D$�$X�@��ų����x�� �"���mA��F�ԅ{�)��O��ȣ�٩;�qzS�����[q�~$�G�{�ĸvh���v�2��/�ŉv��)��G:K/�!���N���b��tժݢ��śJ��,F����b	�L��{+�\N_����5����a�ڍ�� XL���Pz�N~VМq�3���N�ݻ0���w�ܑ�yA�bV����ZU~7�J7�l�Y3��)wm~~���y�&[Z���mp]|��j�ֱ�*��%Uh@qĪ�@2�*�	���4�Nr��V���#�&{w��Qd�4�B�5xL:��f1󝱛��N�6`#����]���N���r1K�.��6��6��퍾��=^��)�L^	�c��1������4Nl��d��t%�/��Ò���,��*�d����5�ó4h�(g�Q��<�?A���t�B���-�z��2��:��<D�<��8���Ɨ>�ZɤH��&�P��m�E�S���l�������m�__��Z�K�"�0r��L�%L:��!�"�c<�2 y�����>�l�E�#��I�.\�ZT��9� ����3�Q�)���j��BЕ^E�J�n��,��_/{�D�E�����K��/l3/R���+k���^n/`���w֕NZ���T�D��Q�ZWw����N�Z�r9!H�T�7Gw��F�۲U�X-D�rf�:e��� �,ay���D�sn�뼥�#��n�h�?�d���M��	/\�G�t���z������DM�z=%R�8��7�W���W^�2�E���D~�5b�*�BbP1 ���Б`�f��I5	U@�k�t�2��Jٚ�H�ꫴ�.La{5KDM�~��/�ƚw���j����D]�K�\�5V��=)ѯ�(���
�&M�t�x�6�%ԋ{�Е�ܣ*��	15�6ot�V*Ie3<����bBM��'�� Pg�?Z]c/M�T&�=��7�#K�Y�"w+�bn�%0[].z��'*�_��ҿ3��̄ph��R谼���`ߎ�7��a0��?B+|c��{�q���y�o�3%����t�L _�p���`tGM�N�]L��_M
��m�t�+�D���%0.8����

Uz-n����#8-bu#b*E�S-\��L�x�9�K?ʟá����6��~�J��C�k��%(��oRA0 �����+�F���>?C
����u�SMH�RSpF���9�$�s"[���7����g��6�4W�� ��,вk��h�VMaP:i~dDՖ��r�[T=��+az���W[a����`Z�0Ζ�wd=��5���{]�Ђ[n�I�i��c���v�6b8n5�b�9Ɇ��P-��G5,�Pޑ`�ď�������!��������G��c$M԰��"Ă������<���u�K`�)�b����)yq�e�e$+AFȫ�0�eM<�V�/T��n���k��7�N���͌ջ�� �F���i�ζ$���i�$)	�s�H5���gx`��ʵ�Ş���B��S�3gd�=��-_T*�o�cz
�E��hP���w�n��=�:��-��*G�N���L���I��T��4�6�h�]��'��H#Y�;a/S�Eq���Φ�� _����ބn��q����>O#��4��7f|��@���>'�h����H`�X�ak0���@:ׯ���x5Y�$�5����	��f�+m�o̹�S�@�pn����n")կ�����{�Ҹ���Dzm4p�0HIa�4������.�MCXŘO�e���=�.m�U[��q���[���Wj���P�ZGC��Bή�T��N�6ԝ�0��#��}s��O��n�;<2�h�4W`hz�סvb��j��:�te
�N�X�v#	��H�%o)Z�`Jׅ�Ѽ�9d�ZQ�*I� ��s�C11�˨0�U(2�62I�|u�N?�p��9�����0�u"��]��Becx+VT��>v��l����M�^���X�zl�w3^Q��Gjg�]#$n�?G�!7Q�ݜ�0 qL!�】�5W�un��1�[_L�mGC��t���Tb�}��f,'zG��3�&S(\�X�V�'0��'Z�z�;<���Qz�M����Ƴ�Ƌի�aZ?���P˿'��� ��Hkq,�`�ggZ��aah�,�-���b�\b��*ˋ|{�j?"��,5�p�v$�҉)�H�u �(��D2��$^�Dt5�����D�c!�E}���R��W�M"�4t1�S��O���Am��7i��7	�ix�DF�V����2,9�*����2gD���NB���@���ong��ÜZ�
"�"JǼI����d�Jr�?����j��ria��'�ߑ,W
���%��$��CB�3��WDڻ� �
�&�f8�h�<�D$E8���x�n�t��S�B��4�L�w>��z`h厮�6�F��HÇ��Z��F��`���yQ�ka#8`�fٱ+z��w$W��`��`�{j^�ۥ�qI� n���ֺ����
,ǳ�����8�1�488&$_I��#W��-�3�AS�ъx�,��@��|����Q�����[�N� �pZh�ϓښ(�(��f{����%^xY�!F»)ڴ���j�.�%,�j}��þ���Fw����W9	�2��Na.�9�A5�IlX��%�Lz��;o���K�%;œ��Y�T�.����Qw�@�S��m�T�<�]L����|\�R�������,U��՜Ϯ��zK�|�5{�$RL
�����Tz�'XUq���ج<r	�*������տ���ft����Э�:��4�w;2��V�.�������MN�O�����?�ޑ����<��<�3]o}�\g��n*P0��p���ɣ�F	^�Ыk(b�}ng�R>������ %��]ޑW�J�r	4ӣ�;vA���q�y�D�?���+��{���/9�$����Ne�٪$�BȢ��GF$�m:��B�kkڈu�o����=P$�g#�z��<m3�S������S����E7���H'eQK�ѝ��_�UE=��e���Ov��h+��e�nܤ�ɩ����H�4�^�Y�����c_zا2�@`[rw%F����S�|��r
���F��4^��f'H���=�2����B�3�Nciِ���I��}��Of*:�P��G�eo�;����p�����i�5�kTB��9��A0W?M5	�Z���% �EW��&W�y5���m��:ҺJTImt�� :����(���G��_�XT(0q��nuן�M鰆�?RX��ǢwK��`U��+:�讥����I�YW����a�@��C�'ˎ��)fT�_���v����(��i6G"K#��!P `?d!��Ho��u*�9{�#�|��������I'�U�܀�|�b4�I�A�ъ���=<��y oBOJ��Mf����n0��Q#|-������!
T�KA�Y�a��%x�P0�IS�:`�@<Ҷ��0*ʡ�%Y�e�`�8��P潩���������ڨl��IѪq(��DIf)xs���m�կ/S#S
O���@yX�h�`E�d\���_�6j
1E�h����� ��w�K<�kr5)y:�ی�"��O�R�Vf����vg֎b�*}�eI`��(n���R���U��,ڇ�s?�I,�"R���k�t[Q��3�l�l���[�����m������Cbl/ݍ#�\�wT��<<rޞ�jW�\|M�n��W�Y#�.(g7�\d�S�@��U�:��i�����K|�[��z�7x�H+�ڂv<�ٌ	-D|��$s� GĊ��~��8Ql��w)����cn�1ei�b�����9�w�yK�f=��و8YBd��mWT��,r!<ޣ��&P��N��Р� ���߭!�p(d��8�h�
s��[Pe�yI��Mݎ��tT��h��}���$,nN��i�)z�)�x���F��C˸�Rl��Q��@�D/��#�I�}�Ŭkd����_��}�]���]c>%��Ua��F!D��^mx��~���W������_�F���>��DAV*U��u�����C�7%Z��$�˕r�{`I����4ڟG(��R����W���Jg��aZ���Ή���֬�.Q\W2�w�9��\A�^��k,�%��<��"��N �e������غ��4�m����OlZ�H�Ȧh)�\�/�����D���\��8��Ob�4�4�t^�t�)�诛iC�A��W�B�z%��j�@VL!�����+�P+���J1�z�zXU�����~��{����bgY�k8��}s~��K�u��Ć��1������oG]9�j�KXr;	�@�����pN}�:S}gR$�>�B��ק���z��L�n���m��"����8�0��/V�.�ު"��̘*�ݐ&W�6�������mJ-@�i{wKf��b���XM�� ��ϋ?}Iaڱ�bXeq�\��b���	Ы�������Y�R��$�տ4��;�W=����[�/��DO�NM����)�2��h��ɒ�׀%�g�M���QԄ�p�zH��_�/�&Ds�3{�i+l$�D��0C>2�S?X�8N_7�(P����z�A�G-�z1ak����qN=K���yKͫvwEe�V��u�z�������� 2��F�A�ن�M3��?.���_XUo(y@r:���N��o|^ _�y㄄ҟ�?N��&7W�>���դ�Mف[�';³"��*E���!Q��10�\�Xw��d6��ٯ�����T�Xt�6�%�Du��O��k�p��F�����H&�=}���EQYw"�K�t�G�@~�6��/N4h�MP�y�@w?wa���{F�̋q�D"J~�.W
%�^��� ������&�ɣG�eJ���z��Ž=�$�#�DT4?x����f��^w1�b��=!�K�9v@ �H�I��TZb���j	˾P}��V�>@�v,���6�����w���-�e�ѢP�;��D���ڴA�����q������J/���=�Ȿ�B:&0Au����E����Y�˝��ky�(7F���6O�"���t�x𣟖g��E!���:{�FH[�8Z�V�^�p�\/o����G����d�w s#0&+��s��]^R.K���r2�����|5��/��@������M���X�j�;2�Ѫyb�V���6��P�ޘ�Qa�0/]�tc1�.�+�\�C����&AhF%4��PWi<��L��R�V]��)�?>�ۮ���d��<%3�;p<N�7R�e�߉}ʬh��;���1Lj���H�~�=O7+W�!N�����8�A�D��%A���/�H�.�(�����͕y�1v��H��z�J�k�E�������'Rt�R</��SVoT���8��'��P9��4�u %���EUĒ׾)���6��?s��]�Z����_��F������H= ]F�Gm��8s`���4r`d��s�q�Tc;&�I[�x�kr����{��wS���%���e7#W����|���>����iK0�&������8@}��t���N�a�j[��2����D�W<ŞW��{V������Z�zj�o�M����/wtx��#{�u'I��A#���h ����KfՇt �{g6ʾ�R�86�#�9U�ڦ����\�]M�l� ����h��gBh��Ae볝3����OQ��ϖD}�_nV��8."�#��5ڄ]�n��y3�e�0
�D�f�+���Ac	��=��I�̒�)Gu6-A�������Mh�o�bG�H!�=I8�&��ǚ���*�7|&�������Dg���?î"ڄ�x�B����2��>9[ȗk#�7T���n}���n>����Eɰ���2h�$�)*0̎�%hj�7-�-[�$�b%2���al5A���h��?���S�R�$���@7(;�~v��e�)�˕�~�}HCx���Z%�@^C�2	��!]�!m�������U���*��M	;���Ș��l�h�:��!�=�6n�-s�Н�{)R�^Z�au]㤯wp�2r�.��';	��[��do�B��=�tT5�EeK��_�����؃�SQ+:!��0m(`a�Az$�%O,A�G�s�H�y#��W���-�Ԅ-�5�,� ��6�DY� �1g�2^�M-��[
,TI��Br�O8�T�V}���~���O��3�r�Z!��e�0�cjY�߮���N�U'D����_�s�En��XHUT��!0R���|�*?:_��c�-$xi���S>���A�ɫ�+k�s��qՎ��)��qե,�*)+���Z;�����w-�-k��3�Cz.	 �1U�<�9AO��5"T�O��A���d�a+������Ƴ$K��9]*���Z��g�;'"�������WHU��ش�̄�؞77����,��Za�d	�:�r�a��H�!d�z�#�fE��"I�'��1`�{ۆb�&�'�;TḊ.c�:��JZ�S���g�&ݽ��*&�oo���x2_����Oξ�g�O�G��=	$��ݜ�r��Pi�,�PNOu�y#�)�'(b���nA��t�[�3�8��T��l�~V=��2����ЁZ(|F�#L��a��3s8g3�O�K���՜I?�0��=*��e��P;=A6����W�K8�%�R��}�J�������"�P�C�*�P�}#Itk#^��)ħ�y���(2�r}�j����W���]u�~�(��DWK�L�L��°�#�d_&f�n@ ���4.p��~8��Q!��"�"����9PV��{���3�?A���'�J���-	�.`0v���[�G$��t�Ī$+�B�R�i	$��3�ߖ4.��"���5�J�{����Ɨ7�E$c�1�4���eË�o���I�)�������O���	A�=�R���5�
��7@�,ZɷoC��{�m�Z?�y��?�h^�wX.�����\���_#X"tP���.�}�0B�|(}��&�t|�,�Q�z�?���K��y��ȍWk��+��4P`ے^�=�E�����ӑu����N��@Y#E3'"� >Ƹ�B�-�hc\)�k
izW�B�$S��H��]#Pa�?d�S+!��LN�������Ԇ�~�;��������䌊-��+h���׌�7�ɿC��ך�LB��N�g����E �g�:A���E�&�_a����eJ[%*Fy���\ �����.�=J̠��]n��nˌ�K�0�T�U�Dds�)-@���#}�Zs����LK/EO�8�
��&�Y:h�w�;H�M�$Oi����3�C���D/��4���AOU�P��I�d� �.#�Hi�K�:ٖk�P#�t!���]�e�H�m �G�BԆ?�E���|������rY
�A���֥5l(-��#�����n��)��/����j�ZX�h�HYc]���v�8��}�D�0�s!B��/K���p/��g��T�Ih�S-mF�oa4��Lp���k���Q�Ԉb߼��f�	�H�{���I�������7q!4琲��펷N@�@�c����^����7�������d��+���1������55">#�D�Z���G���U����s�V��j��e�!�X��8�3��i<u�O�fM��P]ө# L{,N�z��������{
ߊR/����"(�ME$�����C���c��֝�h'r�xz��
jxT{	݂��)�C����)�~'v��e,�� <����C颽ݫ^<���?>��x.��D�w
�(ZN����K�;���B�K�:�t�s�����+��ncd��Zi3�G������{������ʫ��n��͈EU�3�Cp�_0�|���#be�X(�9������A�=��w���1.��s�$��i�omZ��������L �֣Z4)M���ӗ��G�'b�#y�Y���b	oCp�A;�:^�FH�JS��8>����l��2�jq,�J������ֿ1���z���9ފF5O.@I��)�ͬt�/aeǅ��p�4M�(����C��n��W�ۖ}�������Ekv��ׁZ��:N�<�H����4j>��g��>�q2��c�������ib�e���Z�3�@Zӈw�(,�t�RL��n�y
�i�	��τ{n��P�&��^��*���U��*���\���?��8$F��Z�N�Œ�Q|Q��V��x��O���ؼ���XkYh�LL&FE�E��]-�j��Xu*eEp�U~BTX�����Ҁ��ud���>>��K� �q��7I_IO��xb��s�y�8�0��鯰��<�b��"�d���z�Z�" ���K�D4���[�ӯ�
Q�ʻ��I��������-���=&|��IԄ9r��C[t��
9 ��E�a�{�YpR�
Q"P�s����9��m'Ĵ�X� l�n�{�ɪ��@��H ��>�϶��s�r��)�n�d��#���vN��;�^����E�7�urg
B)ujpQ��	���A�߹��������ǔ��r~ԙ���>��a;J��۹>F��� O��m�9\<�.���ٵ���Z0��[�N	�I��c�t���5
�m`�)�Cj� �]�X��B�J��Km���Q��dȬ�'=={����R/U�Ϊ�gq"b�X���޳l���ZX��F�
����~G�BV�­��N�����ǜ����v��r�m!xvR-��\�:���Q���m���y�o��Ǣ��Ǟ�S�$�w�V�i�"QY��Oʢ�!�$s���T���:�j ���~�>�4�D2OwT�i;��S	�����԰-�'�!��)��	R,1 ���]��(T���d��A(/��!9{��f��'e��w���숔8�]xSM5&�k��SOs�CT�	��O0�E&�8�!��i	XhM��s���WnST����&mڤ�7bi	��e:�L R�A�kC3y9�rI��p�b� ȓ�d�J�Ê��Q3i6R�	���]�Lk�C�S����@B�`jm`�9���=�J!������ӓaR��cy��;���
��%�?���ߢ��#�K��EQZ�`�,�3H֎0IY�	�I�Y��.5����p&���y4�E�OH��!���QAZ��bMu&G�~Ə���c�@�,ا��+������"u(���Fg!�GYy�?��b�ph�oN2����8x+��l��ˀw�b��b|R�yB��\�HJ������K���s�g�ZϿ,��6��UV����[!��ŕǿ�HP޶儧���*���i(����U����2�ۃ�D/~Y��f	�mH�=;���:�/f��7�v�S�������݁�E��ؾ��^S�.4?Cd\ۇ芰}�.�w��w�1�Ih�d��(mC>N�;VaR����{�%�f�>�L{o_ȶ���*��]J������p��z�uv���<FY��b2�*�9'�c���ѯF�;8IhNN�?���?aʩ��&�P&jPb;������\�#��-���W�U臱M_��=N;ج�+�|�[G9��.�;����D=��s��\�e
�Z���o�%�����	"�!F��pnu3���ۭ�g���C^�]�X$dok���9�Abr���J��j Á�Ak�g�=�%���q�;w ��~g���#��D���U���K����-��hWop42��C��X�n~���dl�x�bF�(���6��rf��ݺ��t7��6`O�Z�����`]�I!�Q��cKo��YZ�K
��*�#�a����_��8F7�O���ʃ�CJ�Ƃ���cW�.k(n��g%��z},�EE;?�G�e�E=ڝ����3 i��,Kq�]GЦR�̱Tn�/Z�hRt3\e���-=��r~��9D��|/p*���3����m`�����d���a�OŊ��h8�����I�z�8���#:1,�Y9Zb� ��H�Cg.���F{��q\�/@��D��U� ��m��1�S �G_�t\͂�<���a���ԌsU@�n����G�\2�s��G�B�n(������s��~^�+�+��aV���Zk�������L�JMC�:��5']Y�mF�)�?0�9{δ��_��"9	zP#�ݽ�4$=��M�>�
�����~�=��99ػ�4\�=�g��4~�:�*nJ��me2jrB�P��}�/(
��=��SO���3B����&j��]ڦ��{��d1�cǁ`QxW�u@8o2B�a���(}�3}��5������ƈu�T�B j�"��5���n_�ɕ�0�����WH*�%џ��R����,�l��X�%.֒�x��"����u+Ү �21�Vr�ϖ�zd�avhGR(��A<,��(M�3u]{�}�gy��ʲ��i�������vs�$�~F�9[�S��َ.����8����K]&.
�,�y��#���ܵ��+�C���n�6�+��aǼo�9���Lh�sv�54}�}o#J��t.�G�;���T�p��=I9f�Yi�R�L�%�wjf��"���L/Ǫ��l�����;:�2:{2u���?�~ ����x73����L��&�3 ���T��F��|kd���>�|�!�f��ƑC u��E�OC�hXg��:��c���(��w�'XQ���[�A�#8���+V+���( %֐�מ�Au)�'���*>MɚWJ��l<~ڼ8��7s�h����м�~�e�g �Z�Q:�XV,�=���P��>�.�@5�����7�;�~D��bM{D3�Pad=��)%�	}�S7��f�F���w"�zTIv.A�O,L^�π��[�?�(t]1��\��<8R���]0��-5"��.����V�ϲ�`�r����}K�z���\F�� �Ys� �h��(������{׳����u�����8�Tᕐ�e ���q}�=5�"�YNH#ʣ���Q6�"���b<��Yg{�qS�Os�#	�h��g�U㧓��g��F5{������{���S�������ȳ��֦�{�/\�.�aM�����(v?�e���q�=��E <X@�P��6q��!ӎ�ؠ"o�ݢzʬPD����B�W�d֏5�v��h��S����ēAk\���s �Ԅf�;w�c��{�n钊F|�1s_K���b�TQbh��2~�f�	Y�O�<7�ܾ�����.榮<:*�^PP1\ٿ�b����E^��Q
�����[!�'����q��'�>(x�;|��ݱ}k��V��&���7R�;�m�:�R�	�� ��sa�")�Ş/�L*w�����MeV��Gj�e��]xJ����+u�-Mj���pف�߃�	0uX��L|�F�4�'�d�өm�$�E3�uI�����8ݪ��'�Ĵ�<�$r�<ip���0��e�ֱp�D%�yI��0oRWz�Slv��B�������Icަ�E8���5�a%��	N�AEvB���*D�����]#e�v:\�-
	����>�����it�����9{�RdU����y�~>2^T�n՚81nb���h���X$�QQ랅J E���N9^��Nw~d�.�EP���G�)v�ֺl����s��ݐ����/���QY8{���m���槅����?Lg�:�h��
�����k��	C�J�Ӻ�l�7~��y\6��:���;!O	Dx�HM[H�w@"��t���9s�x����M����bxb���ż���/Z�,�ˁ�����"lU��U��ǩy��G����1���3���bY��Z���A[Z�99PQd�<#��.o� IM��Ӑ�M��|�tZ9%���h���,�"���"�-�l�>U����3�8{W~��p��q��E
�����2s|��3��CkM*"��q�R�Uv�d�0�KuQ�"� �i����"��`�[�t ���Z#����wÐC0�lD�݅�&zay��{��,5G��D�\�b��L�����Fz��]���&�����i��'q����ՋQ�1�T��U�@����Z����g������P�'n��|$�&7���Q�Ѣ%|W�/���Y�CSםΒ� ���,���.;��S�$�w���9��N�W��6��!f�UF��H-�%J�g��3�je�c��dى<�����N���5%,���ri�7΁��0�j[K�]�pꍇ�L��Ch�+�H�{k=�n�n��Q~7=��b�(Ew�8q�vic�)�uv����1�g�6���>��!e�%������Lo�<���da���淋?X'�,�9�MC\X5��K@��9:Y���&�`e�C�A&���zC�Khad~
���>f��SJ���Ƀ���X�3��oB��-_~�f!��z�k0�<��;��l��cB�ĺ�Aѐg���'0m��"f���ƨX
����#�Ƃ��LX�ZK��z�
��A����2-#���	K��͵�� ����H�P:�,�5zg�g�iA�kw�������tt�e�4�	[��8��l	��d=�����J�+�Yǥ��Ϛ�\�bP�o*��X�=E�ݯt��"۝�����B��0�1��>�T�K�L1��'�V�s���kg���8��,����o7�-qO6���<6O�a��gu�9j^,p`wIy��o��,Q��\P�|�&�z(%�ҧ���f◍J�GW�k11m���:!cI��񌾵8���-�[���ĂC�|�K~V�`�e.
0~dP�%���6��T��e�I�֫�%i�I�Yd��!�� op�!�����]����������@�3�'�-�J�g?���-�\�3���+9�ԍ���NL�М���<�y���N��l�K��%ôj��&���������qv�`�}�@c7$�dZ�f�����V��������P�G�%Eaӊ�ʂ�[���s����E�X'�5�:-ڤ����^Gs0��An�!��s;�@Iw!v{0�:+#�F���(�ա�<���FԄ/��G(��Hq���5�}�p�� )���kkUQ�/����Z���p`Ǎ��y33�w��?N��msl��?e�� �r��޲�v��G�e�}�o�`%Q?ٹ#"5~1Tpqji9��sM`/����1�+8����N2W��(�������z�Lܔ'�J�n�ި�=@d�O8\٠W�H90�}��YW�ZcLU�)Cђ�;�yrQ%ᨬ��=t+/F�D~������nś�H66sr�����3C�|M,�߹�͓�)C,P[���:�~ �ga����.E�o�TAIxz�n�Z���0��B���k�$g�F�ARd@]�#�V	��OH�;^�76��t>����31���Hn����������)�Sc���z$�F�2�C�䒹M�FL�M�!]� �%ʽw�y�1��9��qI�0b����'�f�dG��Cߎƒ�`JHާ�1.3_/Z��QH��:�L��W9P�l�_��Ke���&���z!�(��.�;������p��A��:f��n;,�B����~���z��)��F_�t�Y?r��ag�"��ݺ,� �g�2䍼͝��UAv�@a�z��UX��1�D0���1T��e.�()
Y����޷5^����|��֓�
h�������l�aq���|�7@�u~�c�Xme5]�����izF"���<xB�u>e��\{y%53AI����dE/�ݠc)w��/p������I2�`��Bҽ����GPt���8J��J�f��7¢p��h�
�z
�$��49�W��ba����=ϖ�S�n�&����8�k���;0i$�9^T��W����̤v�4�e ?*���4vx0;�Qגć{(j��D�`w�L\gQ��H4� q8��p�-g�nC:ʌ%h�u{��͞�R�!��}��@�"M���Gs��Uo>J��A`�2 �u2>g=�8-�S�u��C�M�s�hOb�C+�n>�N.��괟 @�a�¥L�6J�"H�s��x{��4k�4У5B�M���\���T�"���yk�����wc��;�qZ��Q�z+ H68�M�o	^W;j�\�=��Z�M��W⊑�5TGLm�w�:�`����o�4���R����]/�Z*|����%C��UM����,�le.K���H����~��J�d�]j��v�PJU�����_l��� ���l���<Ϩ�a%�����u��	+�K��2ku=Dw��Z�;6��L��BJ[�X��F��	a4M]��Ŝ6�؅�`W� ��m��5 �� B0X��6�JI����_/,e� f�/�6M� J����i��;�K��4p�� �E�V��t�k�L��Lg�>�m.o�.ԓ���d��~�/��W|�k���A���)B�o�ft�*-U��>�p���ݭv�R:�������<�"m�D�v3����至n[��	?}E0moMt�A�q��"UW-�l��� �6�q��6T/n�f
N�|������4�����>p�|
$�)$r��g�N�,	�(è(�wZʌ]�=z���@�W$ 6�n��Ma�1�����Dk�S��ȬL�Cݳ暕7O<,]�#�U��b����wV�y�Y<�w�s�l�Tv,���|il�ݙR�w�%�k!?Y\(��ǉpuZ�je��͌��kA��О<c��m�-c���@%�P����g${T�F'*�Z��q���ƣ=����lK]���z��������тZ�7 ���N�47D�Ψ�⏧�
#�{t6�
�o����F�o�Â�����p�*�m����5
��E�ۖ+?O�m�aG
}b
y��8«�2Uo���� �<7w��uJo�;S�#�_���x��5<;˩@ ��8ǐg��	��i#)kk˶g(��>��/��R_V��pV�|�D�Y�ϻZf���jptS	�2���=OBm�ʡM�9	OY%�a�QK��?�
�̢��F�*YV}������<fu$o�H��~�ӽճ�؂ ��	��iժz���R+]ۊՐ�T�hM���lЬ �$c��ԑ�]��ʑ
����D����)�J@�t��H7I��#�g&3���Hl��#�,�����r$�!�p���n���L0ݲd�ӫ��b%/H�8oǭ���D������}5�u^}�KeM2G�^c�q��,�1�`�tN��\�p�g����p��S׆~�o@u�r�@f�.�ڬ N��/Y��҄v�zr5s�y�&v����p@��L�)}��)�¬o�O���2�x#_�+�vEPv����{P��>�3+���Ro#Ղ�@�}0�g�ߟ��mӫ�hp�(�0�������)��>�	��d)��BI���;�a��,�Qu��b�Z�Q�V3�{ ��#��ݺ�вS���:d��|n�=���+�V����<��?���Ԉ�h5�Plݽ� �F��k�'�eo�[v��IBA�27�\#�V"}�,^�E�@*�B�$E~z�����Q{�HYe�I2���$���N4�����1s��L�����AR�����?���Pj��s��'��X�y)���l���X�;�<��$=�^g��*��^@2�7�ݕ�୨�Ŏҹ9�t}��z��f����ٷ�_�i�r��V�O�|��S�n%N��T2�^,xl���E @�hk\�P�f�|�oV�9��L���E���by��^/�,�1x���"39:�AU�F��u�ڬ=>�݃�Y
g2A�4+�1�F6D��`tN.B�CZj����WوFtV�M�C�H���kAG녤��RƷ�J��̶>�І���30�J�]�������<��h�����Z�nSȇ��d>�(�+0���R�C�=�jB�Q�-��	���c�'�t.-���i�4#��'��kV�$b03��،���z�a��{��O����D�w,��ok�h��Z��{�>�Ğh)��-����>C�{1��q�\����26��~j4�[D��(�{�?��F�2l�i �����;������:�̸Sފ'���H��WH�W���(~�^�ƚ?����1� �ݻ�\ ���F�g�sw󭲣�'.+�<'`��~ht��g�P�8g#��o���vI��\�%b�HB>;h34M� ��˝]]-6��aH�}��b�9��۾�!(��i[�x@^H\8��0�a��(�v�TU-b��>� {=.��1�G3Z'�+X��2�M�J�P�����Z����94")ڇ��@cv@89�<�g���NFf��� �$K�
�`itBm�t�$K
-�K�L/����~��4�fB��D�|��f:�v����n�.ֹ)I��:���t}o�8��[P?i-�@�����E���B餸�O.�v���8ٔ<:�7!o�v�����B�m'��y@Q��g�E8h��3�(W�`�wWax�Y��T�N�\B�]��N/4CC��W��;�1����y�P��v,��%Pżt�?��Պ����v�� c���fKm�^}�Qeg/@���4@K���iV����%D�2U��$�^^�&튨-�e��$d/�MOÉ �2��mǪ���M��p��7�>el[�ᦿY-⥠��-~{�Z�P��fF��gl*E��i��3pF1��X�E�)���q���A���6���c���ܙ�:I@���>zg���]dP��L�@��\���q��m�&d�����,�2�5p�����7B0Qv�;�w#����yI�*H- T-Tմ�7X�ludսz��"\��գ(f�=��4����z��t%X�y5�XIHg�
�y`m�`��{���1�_y�ʝL� 0�d�����i��K�ᬲ���'�Y�:2/�����'�
s4�I�n8J5�8�H���ze�w�9Γ;�B�~p�~�Z)����zD���ʎ D���n(�b$$��5���]�!B�t%�3��y�j��r��/p�D`�_>��K���FNk��� ��W�g�~jW�M�z��`̼8�Y��w<�غX�r����"؇�����g}�s��Ab�E�:�-6�� c��/�B,D��,��[㠱w�<, y��/A�{�����O���c���~W�D��4�d��P��d:X�I�R�93�6h�aL�l]���3ܾ��}=��*���G������i٧,�{Ӵ��t�i7�c{*~�O0
��FѾ�G
�����8�;���']�8q#ݫ���@h��Nķ:М"����{O�=��f�w�̈́��'�dJ�	�q[]�9 ��IT>N ܆�D�ŀ���O�'>`�KL�w�����Nᆪ�.J��co�'��	u^,��"���N<Q>_��~�N�V��5K�N\�jT�BQ��%�e>s'uv����+�q�#��$��_�V��ܶQ$t�}�?�56>)���6���iS�g�NB�ig�� ����l�%�WѮ(L��ޣ��8
{zw���{�s�l�f�,n<��uw)�!�z#��݄�>�~�:����5��!re����IMSB��:ڴK�T�1�ܚ]Dɸ�R����wf�#u�o��[�v�}}%��m��[Pc�?i�L`��)�J�b4 z�����'@�~_�U<Z�m���wQ�9��g�.��*�`o�<��oE���_�|]q� �`�x�*��/���tF�Wâ@�<�r����`���	"�[%bʐ���v�T+Ěyj��9�n_� ֯��?�nAj�R�|�s��lr�5�$�mY��D\�y��H�8U ^��dJ������nQE�W��
i��·��y���D�4�3ҿ�s�Ȅ�œa�^����#H��D�O]�3]�b۩�c�S�IpI�J='Z����MD���7
<�uF�C�QM0K��R�s������nK��/(��`l������KJ�N�#_����q���QO������2ͧcx��]��׀�fټh�_&�`jZ�4c!��[�%�C]�	�苈���&%�2��)]n�?�c��.�-ח�n@�����؁���dӯ�#�Zvz�}F�!��w/��9m�|H�S_�-:�V�v��P�yx{�i����q>��R�x*R?Y�L����/kt|��/R>�vK�V���S��=p��5��^7���h�S?���3��{iBi]f���[�VH�ZT	���X�ٖ��ۧ�s��l����\"�_�p�w��c�[�M*/������8ա�{']�l�{`=�����6pX��m�_�p'���Z`Q�O��R?Ո騤���IG�2
�t�;�N|t'f3Y;O����Ʈ�X�����4aZ��z��3G�a�˴�se!�!Mf���s��5)��V�R���_
��`ퟨZ��FVβ��<(X5�L4�/��#R]�4Q���G[뒠B�ec�"�~j��J����O��0p��|o��F�]��f�& �NuI$Ѐ����.�΋CRWb[j��p�v8g�L[F�h����O:�|��?�ef�{�^0p�w)$���7���^)����)�����c���J}I�=�|�(\uq�k�Q�|"(p�~c|��S{zA��O��
��ڄ<��\Z��	�䃑�˷��ܶ���c�����v=���V�̊ߘ$y���k^��`N����)1>IQu�oP�`�<�sfچN��[�/��t��Q��]+pm�Ʌ��}����w�b�c�6� �0g�G�s�/[#K�s-�V\���<p��O�9��<fw�ljQ�u�7�_��)�br�/��Q�^)W�qx0r�<������$���^u��J�+TK&(�h�Z����K���6*]�,�i��,���3]�8-z�%��P�"�}�""�=��x)�D����ux�7�9�5����@��Y�Y��cf?��U,���0_P�t\�ifdG%�Yܵ=XjE�\ś��\�O(���,�-C^l?;�؜$��N�\����Y&���� v���BnB��>�	�!#�_O�Qu"u�\�!������b�� ��!��@n�M�"I(��{�֯T�C�c����l'�Z��q��ۧɥ�z�ָQS�oQ����&��sT���T\j�6�-�y�6�c24��j�{��q'۹�T�$xYn5	���x���Q��p��wr�FX���܄�RH�S��!۠L��J��=4"3,�H�Z�X��CN>R���b#��dK�2|�ZBO�|-�^�r���b�Dk��,��ts�EM8@4|�-��8g|:v�-�Zj�B�R�0+�]��0d���DnWʰ�e��ҹ@�+zeh�P����]�����`C~�x��PM62�@�ǉ���:�w�]�+1��^�*h�q4�5���{�,33E�suc�1@j[(�+�{�y�.ؑ�'"	�H�����&WoE��h���)&�à*\l��I�ik��=x.����	�Q_��g|,j��$�v���i���ŀ����l%�*\���xi�1��&�b�G6/5���N��&��'�IԤ��o>��'-o&� -w{�i:�[�K�*�4EMw�o�'g"��c�C��*6���Ȟ��T��"�3��,�����![�Lg�u$e�'���\5\�_|{SI�}��3Gv�:_�d�9��V,�L���v��X@�ό� ֱ+$��H�p\��	fG�qF�K���J�
�+!��ɝ�'�2N�,ۜ���?��U���tr���8�[\�����g�1���w����q���>N|~���Ȣ�Z��X�Io��Å��'�3����Z�O�/���|�O���:U��J�����ۇ2�&v�Ǯ����1#��t�a�D����G�8m���Np0����a���x�
E�v[;q�q��p�mv����Ӌ��&����燊~G�Wݑ<����D2���E&:U�1bт�w^�eI���1����,�7DB-Bˌ<	Z�������.B�N���x�y��Uז�٬�,�wǬ	������sY� ���-���.�B�~R�gJ���x�)̭iu=��ŗ��

sk!y��_�75��>c<kdS�ڒc��ч�$��_-����|�R�jA�Pdr&?�=>N�p�k�a������	'>�����ɶvc������?�쑶�7R}��x,��@c�M��غ4W�� GSF�P6Bu:���W@��b��Mё�"�# ˯:[�p�FC^���!�R�`o�d�Ob����/C���h�6F��ӿ������Y2[�Dq61�~%L֪�lx�b�x��V
���������#
�i~p�w�,�~e�!���p+W6z6����`,�J��+�	�\�׌o�vJ�v�9A]E���z'�'�Y���p�)ԍ_&vS	��J�����5���޹V�o0�2܀���@�@�%�Q�Z�l^k>8����0��B�t�6{ �~Df���0�? )}.?�u�"� W�֜�_�����Y� �P�4�8�)+&ZL��.�oaS����ΑHOJ�s�|h���`�hY��0i�D�fGTt�v��"�O��l���_�����HaS%P,���S\A��h��B/Y���>������$ν���Ş����Q��;a%b��s:�mmX�'���0�d.����kQER糲kѩ����і[�2��K\�-?j����`����40c���r.���r��6LE�z	!p�r�f\����j<|�E�Ƅ�uS�?�|>�	��
�*��s*�z~����x?���I���#��R�a��2�:�����H��鈴nX�c�l����*�|���1\��R�{�,��şm΢I�!0��il��D)��DF/�u=o�@�,�5Ҵ��������V�*���䭰�I�XJ�F���bp�����5���R��J*M­i2<�� ��_RE��`f�`����wP=C���gY�����l��\沋�����t���#3�Q��p�tK��$w⶧��.��^�n���-c��O�]��t&Q����q�;m��n�S����,��>ilN����O������l��[
C*r�N~7B�bC�'����j��d��[@5���(S�v��:_���V�2o���F��8�D�� ;�V��I�)d�S��h��ֱU�1�Y<���^��*����	��I�R�@��3�f��zY�X�J$q�Ŗ�H�����L�����b�yW�����8��g!5O�����Ql�!��]v���z���Ч^Z*�ɬ����|�+��q}7�8�	_p�'ZS/h� C�֢'/S�ف$�H�t!o�'Ҷy��HaS�"l.W���o����ܶ�D�!�MF����t��*��GU#r9yȮ��*�3ǵ�G�jVk$(�F����M�(",3!��x�vl
E����ʀ�>f9<���"�'"���oFf�����iC���؆r�b���4I�[w�n	�P�fc�����+�Pz4܃l��(1n#��0��c�QѬn���F,Xe�o�����ذHV� \h�4�)J�t����D���1���l}�Y�`L!v��s"��g2?��p�%y�g#q>�#;�~!.sc����ݠ�3��e������;BCC�JY,}5d��۵7Y!J��J;��,��.О��Ӻ���<:W����S��0��{�'_N�߯�W{����a��*�h�m��M;"��ʶѪ���]�ll��7g,�۬$n�i��H-���������|�`A�w/��'9j`�Ԙua>����e�Zp�H@�:�[�E����?��eh#M��V�|�T�Z_2%'m���Sf�%#TS� �a�V-,���,�7a��LN��5��
@`��,��_��H\��E�fԱ,�<�I'u�qo��
Fv~�o��\5&W��e0����[�=����&�&�����^`q��s#��{q:j��-Ϳr$��i�[�Rw�\`v��ލa5��~��f$��v��R⥡䬠ޒ{���d�,�yb9�E�^|� ]�L�	�#�с����z*L��C�c���n��~d�>\w�eq�ckE��N��%:̽�[�� U��x!G�ao.(2�S�Fj��������]a	V8(�wSq	&��Qq$����8��CX�kʍ��	��z�ް��ʣ���� zF�m$p2�?�
�҄4�=SS�c����b�v�����OĜߔ��y\bIq��9�J�d�PZQ��<�����|��n�ۧI�����4�n�=T^�û]��$�[���,y���z?"����r��En59�0R?ۯ���a�����_!��NA��<�Y^g�:� ��ы}a�J33S�en����"N=yzh��?�wͰ��q�)�Qq�: .ѷ���;CՏ�e:�=����n+x�}��*�O5�Fc�ѪS�J�븇���S$ҩ�D)O�/T�ג�yѬE��̲�W���Ғ?�?���B����5�gqx�_mT�i^���{?�i��rQ��X��8ABR&;�C����6A�	�.��<�=�/�j{ta{�2��(K'h7z����V�*�O�>}���<���e,��yG�����%��,Ru�u���8h��]�9-�bst^O>�r�
���xa���Q�������!<����1��Z8��J� ��>��SM8&~�`s0��w������&-W�[ȓuq��o!Ky�j�Y8mӒ/l[YN;���?��5�l6I�}be3�
���`
"k-��)�-�X��4T��>Rk�#4C=���u� 4u�-0��nc��L���,����z�:�f(��Tz�����q�E�`4�b9���6Q������^y��nQN�D�N��n�"D\gv�J5�5��-���0eb��+���AT��o'���4[O�)3�`�]�?1����N�}��˪B�ߨ���"m�q��]I�@;bl�FC�Xg�{+������.N��t�PO~;��B�>��Y0�G�Qc��p�#��ZÕ�eV26iL%h� p�+X���$]
,m�t��BLS��R&Y������b���K\��:������9D����9��pZc��D*{�P���Z�r#�9�&�Y�&C�ؿ�"1��:@�e3	oǛ-F(E*��s�����Ϟ�@P5rjz��(��M��'�3��C�� �2�d��E�Q�D�Oa�jY��Ev/K�ˊXj����&kH���S�+*L)ߡ�>�ց�!a���/s`$/�-T���U���q��+�qF�����'"����XM4Q�>�ݫ�������2W��Dx�y�`��$����m�=���?jUM�Kb8j����y:��$]ʚ��Z3Yш��_��,u7���nm����m�+��+ũ-�:����%:DP��~�)N-@]�%�%�<�6ܕ���p����A��Q�R�R�b�}����f�*?n��wN��*'����/v�V�#t�)���4?MZ�ѿ�c����eâ8r���B�xlc��k�3�"�4<�R���m2C��V�8 1-�L!XӸ7��`<�����B�z�{^������R�[8��-�=�2�DxP[�S��W���`�Zu�A.�}����z$
ďa�3u~��
�R0�3�k���{���$�Y3���ʡp�<};Z1�h:ӱ����EYKr�=^�ŗA��zS��	I���'�N褹T���C��U�<RM/UN���>�!FJ�wzv����ݨ_k4(m"�Ҩ$�H��wi�ؑ=7�ȩq�n5������
�%�"��-ܘZX!f��,P/Xp0��oYҲ�d9b��Y�$�U�l(��/���l\�5�5��,��~^;G��q\�W�]x�ܣ�|ͻ��O����I�,�^u=��P��p�5oh_��aBA�����=cJ��3`�{��-�=�n	`'��P���oؖ���r'|���0�nd�}��P�[�3����ћqU��'Q5�K%ȱ���h�:y��ʚ��D�E����܃_`��� Uu�0Am��3����^
v6��Z��&
�ۘ�]ayb�����GR#�
��E��y�0���V�E6�(׌[b�M�ٽ��X�7f1�<��8W�, n�*�%MO*�QOji��eaچ����q��6���y.�G6�G�J	U��1� ���lU�>�v�۬�����;e��ȹf���z}_������lu����E9y�k�Ib$�F	I�� �H��~LB�4Ɲ���>��	�~;�������|��V�|8�е�Aq���<M~a} >�b
	#ˏ��.L%(]�cp�h���A�㈋HeVῑ���Dc'����qL&���8�%O��Ʌg��<y1��A�<�j��
�']&{aZ��w��|�ףx3������	0p��_�my�@*�g�}��m���;��E���Fʦ��$����:%[��H��L��5���+Q^�Mj�}�)E���2�0C:%Xጲ�SB:���Jٸ33��<��/��׋�~Et�'�R&���ګ���L��;!Y�S��y�R=��F��8�E#=$.�(��LQu��2ⳓ"���B�o�B��(ny���D�KN rk�g�<dP���C¸�A/K߽3i�<x�2������1���ͬ� 9�U[�$�� 1?�t
U���<+>:��p�s�Sz�k��71�\�ϛ\H<����y�Oa׼T���W��x���EV.z�-�����6~��f����#��v�L�+<�#�����+��Ʃ�p	�Ҿ@g�L��^#��}�M��6.�L�4�;������ņ�O�۲���x���f#�ds������T��1i�0Fg԰zJO�7A��a�9Y��/O��]~7�k4��?�)0԰ ��('�Ij;d`쳛�@��������?I}F�b���槮�/��$�d�kM���3 n���jt��c�~".��Dv�2��Ok�j���5��z ��R�Km�.�w�T�����?ޞm<�C �q�l�v\�F?���(eIY-�I�]��*-|yt'�e���2���Բ�+��Ͻ����Fw���Vg��ǯ�ZÐnr��L���jn5)��OC�n|�2f�9]�1QD�s��#�ʝ#��g��L0�v`���R�`���dc@yV0��I)�!��|����[*һ�>?��?�1�w{�h�*!�V��ت��s�K�>�ݘ�%�'�%I÷��u�!F9��p����p��/�L*U������(�ú����[���)ݭ�.V�Q��9�[Y5�z�K/f�8��Ƴ��D�9�"�hn6��:�|� V�$Ռs�њH5�`�~_�s @����!�<��s��d��#Ҥy^�'��s߾3�_� �?g���x�)�À���kt �H@j@�}<�Ը.�����\C+0�f#%rI�|DS�z�[�U� 
q.�Z�1�J�<�ߨ�S@(���I��A�{H��¤v�8mﺝ�Nl�y�K�mE�oy��"rNT��EI9��p�p}������F�t_����P�e�I�ęx<��,�������y�������?�3y@�W�7�F�E!~=a<�-$d�«����co����"h�t�[�d�����O�J� ��}������:M�8��� ���烄!a�^}'�� ��U�m��*�6�?�h�_: 4��~?����@���D�
�8@�GWn�wE�f)V�կ9"��x)�h�UL��umϘ���cwe{i�]���W	��,�WQK1V�,LI�m��[���c�r��|݆I]H���	�[+?Iq�2�:I����e{#0J#a %�8�}.f�����R܌��87^�r�����ő[%x��|�R��3�D�O֨�i�h} >h���
�5�H�Fa�i�����Fe�vq;�4��N�l�V��˩f��p54���viN1KG�������D�^O��U<RS��c�˨o�Ȓ(��Q���aG\:�J�e�N��� �/�b�]�Ԅa�Sn�۱�ӂ��gNg���i��W�5a�n�6�2Ǒ_�#��V�	�22�����,�p���2��^��[�j�f�
�����32�혼� ����=����h�P������H�P��Ks�!ziBPRo@ޏEs9�L)����{u�X��/n��A�����T�g'D�ߛ��g��ce�)�a$f'�,c��R����$,:H�8+b���Q��k?L�ks�ԛ�,'�`U�JIhN���M�S=Ҝ�_[`D4�k� ���Ԃ	���=rgT����JT�t�ĸ:�w�[S�'_�1���dn��рM���Qv�/�a<c���F{��Y�i�r_���Ѝ�&1�I[4,�Z��7_���kJL����-��u¨�ޗ�=���$0x7��G9V_�W�XC? ����ˠ�8c�^q�<�y|S��<.T@" �c�޿ً�`��^���u^���8��}��m��� ,����~d�դ#Ӱ��s��uw��r}����B�݋��<5�)ɞ�1[�Kb|��]<�Q�9�g�.�=MNr���\�'�d �p��PiBBlg\���4��T��5�Ѐ�i2�A?�w/�/�f���Q��s��kRt���F�1�.�>=����A2f�;�
���^�)���cyN]��<�-��/�����>-Fl���!�2�C�}�3O��-P=���Y`�D�.X<����t��5"R�i�}�ዡ��.�4�h,��@��tv�-^/�Ϋ ��o�5,^d�G�EK�~���A��)����Z]�`W�Us�5'�B�\�'��,��'��k$�u�"[�����v9LZeDjbK6�p�M���8��c�q'k�mB���_���ggH�'|�/#w`��h���gw!-B�i��t^��m^d�d�9��w��hz���8�}�jy�1��k�ٚ`�=�݉=���M�C�g":�蒭�ea}�d�NvgU���VE�e f� u�P�b+�Wb��Oɥ����1���W
��FI�p�_'c������Z�ne�����6Y^��z��������/���,�'��q�a|���vQ�&�<t�ƹ2������9xϼ�$������#iծ{g�~��z,+-��u+����S��q�`����wf	����9��3�\��u������6����O�q$@�㷂(�)1c�O�X�4��4��:B�,�fEö;iݾ��XBpⰋ 3�R;�Ocy�HBLɦ���lD�����g�Zad�����T�R?���^:l%{����S=_��k �h � w���ĕ��˲�2(84�Os�~��̜��IFV�[rBA-g3cL�:��Z��Ͽ(s�sܯU��ru@��gg�ƈ	}���>�ȴ��&��.��n�bX���Jx!����f��B2Պ��8Z S?�ERF�iK�����|�H��d��स��%�T:Ht�����a�Ck\�����ii�ˌ��nT��$:�^ֆ�����Ͽ|�Nxt>�\c�F@&u�KJn�a�L:�ά=�h27oF�P�=��G׷ú"hH��6�>w����-&y�;�i8z��$t��z�1|�W#�G�{��VR��%.�k".KaP���A�t��`�y�#�7F��U����moLx]�����tu��5�z��oOen�'�I�;��~K��`�1��a_$k��6xQ΀G���M���9�)צl�H����mT��
�{te���:}��G`;8�R�T�Ӱ�7RS�1�A��=�mh	�@�}���޼mU�#��n���0��bS,��㗲��#-�̔�7ۙvB�n�l3�|��wg�,k5J�=��h"��Jd�^�v�A~�ĥ]�S�o�Yޤ�Y�O���w�K� �ѳ�l�E�"�x�Q�m	�$�l�C�",���R��.�[�сUG�Q��.�TE3E��ּ4B��Ux^�HƢ�ҧ(:t1X3��l٬x�ɳl\����ԣ�;��S4}�\��m�/��jb���ciZ�]����ɏƗ�k.��>�Jq��{GW��ˏ�Db�"D5��M�E�s�lq���B}���{NW��n{j�(��s����F1�W| �L���)]�6�	�i�"W��6�d���A��%ǇO�E��0�ͮNl"`�R�_d@���T%&�>���X�$��|�v<+'�ȩ���L��.����BAB��䖒�z|o~G�vI)�5��_z��Ǯ�ۖ=�4H�K+^	��I&�PKj�X�4<��b�Es����������i}HhFL�V�Slʮ��|
��gq�	$٧ԇvӐ����@�aS�~ܹ�p�
��P��%��9h�ݗQ��o�x�a!��#���s�k�W�R���_�6fg�
馊��P0�@�Ի�����Ŧ��X{h�.���}��*^t��'T���[LEzy���uwT������av8��v�N��!s�3��U5	I�6���*Mx[hYX'g��.L���7�E�h��gڇ�����JqF�?�Z��ײ|��b�/,(X&%}�5!M5_�]fRr���`�b�����\j��?c�=z��<���Q�So�ہ<hx����NV�t;�2q��Ïy{PA��1��"}��)��/���H ߰�jsR�&��H�ڨ�f���]����t-�����$wfE�����.�o0)�q\��I�����<w��_�g����2��un�.�pj?B*�$���Q�0�/6�*Ǡ�d<l�<&7�|	�r�w?��NMǰB���N%j�	#��(���i~K,�\ų)J�A,
/X��{ yj<.��4d!m�មJD�qbfh��w��KQI)���1  ��l�� �Q ���B�OL��9�Ӻ!����:��ɢr`�w�B��|-���y��{�ء�ЩPA�i�Rdn�{ɓT�$Y�P9Ē����cW���P�
�3* ��� �W�+%{i=4D�z�����I{�8/<��F�D���n�{����N5����M��_�˯��<"%��^���/�
"*��	�H�8j�M��H���[�jOF�(����!l
��gU �D�X�����Oz^����u���.��IS��Q,O%G�N�V��z��o��z���R���}RȺ���F2=��dG�ޜ�-@�+���ZO$�����h��-���}/r���2Vμ���:��3�0[�1'�Ū��s��mVP ���e�ד��o	��R
��%/��YV@�^�p{)�#.F9u19;R{^�4��JL��=�a�����{)3H�=f�L��m �uܰ�̚딬;��R�K����.�.�	�MѨ���sZ\gz��ڸ�K'ͨ��P�ײ[Qb�#v �0�9.��/�Z��(q�"h̿�qf;S>hSH+���i�=��uO/H�{I��[dG�����u'��.J�NW@Õڛ
h'�	�v)�
��@�����ڥ�f�eY!��/�p�*����K_�c{��{��B	�S�5��v��������l�:i'X*bgl�NW���X�4����4��e];��6�U�Ev�+�	a���߫�3>Zt��a�")m�Np�=��1�s�;���@a`�i�a��
Jާ��(,jg��?N��*�xK�����a�b����'�5���F�b���w�<�os�ȌA.�Z�Q6)��@M���|B\x�W{����q����ֱ��~��A����^�Xa�;,�H)�Q����5�[��M�Q�CT��	���u@�f���&����C��h͛v��96�²���r����^["Z��e��Y�k��`�G�Ǧ�,#?�!_eK�Bs�@�ʑ^�;�YI��k�+¾��������d���p��,K�}��M��V�>��q)����p#_���/��Z��ת�MMCz�B2�[O��U
�C�;�$N�ʰ'Ԏe2G[=h@��]�{ч�f��cb��G(��1;ݴ�daNO��7���r"8�#~z�1{���]=B�@�������j��J����BښGOM����ǖ]Së�L�	@'�5fzq�21�.x>_9��۹�_r5$��t���O�W����O5�84��d��*��:@	n�p, ��Tb%���D����3�s,Į���x�2|#��@y��cn��s��V���C2YH��7����"�ц����eGOٷG���A���}�.��P�-���l�.�P�
��]*	�=�v�Q��$S��yp�#K���FmƑA,�ɮ�0�36^�i��n��B[���+f��0LUK_�p�u��ϬJ//��F����ykaf��cB��������H=,�ǝ��r��*RY���{��P.����j��0[dP9�����_Y�}�����|60=�?� �L�3[Rp�P��"	8�7��!�IJ\ڟ6;�C��jӦ�*���> �+�I��W�W�G���6}� ���54�
K�m��zb�X�4&�}B��=Uߩ��$��5Q��}\qU� ٮ���#�$�h2��=��d ����>a;��fźϥg��
�rJ�j���Y��\���E�X\:�.��e%��J�Po�!uS��Lqq[Rn'�H����M?ӈU	7�ט�4:8ʴe�U��� ���\`��ʩ��ݫ���=��:�=���
P�8�>�w��b�	�*�RSzt�ģK��7�J�v�U �yJe�fe1�+�#�c�b1���9�`�N����δ��U�(&2��9di�2��C7,C<��E��5 ���\3�!XvN&��=��'���Z�SJ�sM�)nm5��=�r��+%�my��1��!z�rؿ�ʍ�N�D{�\}݈m)Ar�m<�)^��4_&)�B�{��nM������y�}�J�W�ҷ�<�m3���vR�Wߤ F�-!rnNd���>�I�
���aVD�zx���1�::a����jH�ʄ7�U1����l�ӝ8�z`n�j3+ݡ�X�����4.�F�0�	s�o#���.�3^�7d���i.{�� K@�u�'�TjC���̓����%c� ޴i^����H�>@p4�Ä�x $��!�0����'Od#oe�N,]�H�˦���H���,10�5�uT��/Zu��J�W3
^4~�4\�*��*zo[]T>�::�I����#����'o<�8t������lw���.ؗ�"f>� �`J��1?rV�_����d�7������z��J��)Q̭b��%�[u[���T����7�h"��#�B"�/��|���$ʬg-�������r2��Xü��"��_��N��:ï��0+ȏe�zE� ql'��-q@K0��yO j���DЉ�A9�dy�7��η�Bxr�|�S�鎉��ϵl��j_H��"�bWTH���i�(����E��x��XF�^�'\����Y�:�3���د�����7��!_�+l���u���c/Ni�0ϊ���Z(��QS|JN�¨��YZ&�
��������mցt�-�+ ���y��p�ԋ8�ձ����0��� �8S�!��<8y�w���)'U����-�q�Z�ͳ�{p���ao>��Q�M����O����j�婹1��1�Mu-4/�pBJ8����{�d.Uy�D5�3?��wהx�����}���{�a/��v�׭���W�$	A<Q+��D��jBq���[O�Lf�/�@s�G�Iz��Ի+�~���]Ћ"N�����O���T��qi�����~���u��secv�j%rg>߇���'����p�@��uo�ӭ�j.�.���Vٔp���]�������<ұ6����W��޼��=���xzms��4��Q4V㹪R����=y��K) j��q/�	���>�(�dtV4��oA�p������E�����9D:sBO&5)��X�u,r����"�����W��Sܠ�ݗ�qe�����Y��IO��+@�ڲ�<?�9�an�Q�����ŋ��m相���_I�3R6����Mf?�i�\��Ȓ����~�
�����}~/&��
�ҋ�����#����Rm`"���|{��*�6�f��L�ԅ���9rY#���X$p�<�v�zMP����K��ד#߸ef��/f�����g�����X��:$�~��L���HӢ~�	x���w�P%Zf"�|�Ǿ�+���$��6��)�%�-Q���pˡ_�d�PZ���)����z8���<��2�N�rIF����|��ݼװ���;΁� zuN�v�x�S�O]�˷3͓�ve�muT�T��G��gH���TF�u���hӟ�����&3����tKK���J	�	O>����]�k+!|O���?vc	j�<^���&gr�an�Sfv�u˭�4E���8��c@�K��նGPw�V�E�3��ݪ��e.AEM�� �:�
�4�Y^��o`��s���#~g�gAb�Ȧk?�1�����ćy�X\}��0����.N�&�֭y�!m�qX��=��g�(5� �2?�3�`h8�x"*��f��J������|�Բ-�D�,?��(��e��e�1�YZ�dq�e"( "��LHa��_��^pj����XB8Z��gY�~j��S�]�Z��&	"KKˈ�i��m��t��Q�)�����x9Ҭ�d1�O���.;T��$�nbq+��#�{R���m�1��sk�?��M�7��ڣ(m+���Î�%������z���_��^%@�o
	y�i�e��&���b(!��7����?�WA{���%[=��ĀE�ݎ�-����.�j^`�&*�n�"E������l�ia���S�.�#����ہ�D-������s�PT�RAKrsԎ����)]B��N��7�{�K�[v���}p�vq�kӮր��YW~o���[,���tS��}�����]��='��ՠ���jw��К���Z���i����W�(��O:���=a�H.�p� �N�Ohw�|�o-R�Yw"��<9r�/I=�P�� ���I~&Hs"ؚ.�ó�ז�#����)$���Ka(���аS�DF0:���{ir�=���:^�zm�(?����8I���hk+��g :��^���R���@h^�D�YH`�\��m�n�y ;��gw���m�d�*��m7	`�~]ሗ	�+����b�)cP�0�K�)�^��/;���EY��Gf��e�J3�<"s4c�F�]��-	�֥� �Aςe��:H���6+��?��z�?��B�����Ӱw�IiB)A�'2��lY:7�Q�� � ��]��죈�1
_���+� L&�L���Qtտ��<p3ܷ��II�#��X%��g�]�Q(a�6K]_�94��������1��AEn�!Ye�o��4��B4K`�51�'���#)o��H,$l�
���Asy����2'7��
��݋B�'I�F��)���.���Ѥ�}�)	���{8bϝ6���C�%��Aб�p�%D8����M��Q������h���1��a���;��4�����yN��I��|Ba7x�\�OD����i�y��W�u#���q�׈��|���]KPݯ{�3���QRyB��A|�L,TGaբ®���h��"�շA�[�^)I瓯{]�Ϫ��$E'T��ĺ�D�U���V��:tKe�����Qhlz4o��{3��*�lv`X�3�s�9Lu���7���Ps<|�O�1���̭��H�4u�¹���IQq�~��4So���\�h���j�����"#�FV��Q;���"��(�����#=���rl���ύ�j/!��k���@;Fs4W'�wu��6�懅��+w�d��{���*QǩԵ�����D�M��'J��Dc�*��B�DbF9��ޫ�g\���/F�NW�Y?/L���ʓ���B���%������Ò/�Ծ+ј�"'wo�I��{hEsO&1�8���i���e��+Cy�m�
�4��k�w�g�)�(��w1�yj�ŴC �[���4)5*�5��6���zv[�c��5����7�?�S4��f�A�{'[s˽=�Dvli`�~c2+��2ɀ椓"Mfs˝�fҧ���B�]��c��d]��8,S�W}I(<�x+�f�n\��^�Y��z.��GOB�v��R}�<��ⳃ�V]�<v�;������Z�l��,� ����hL�:��V،�C;� -��Ť���h��i㦒�rw-	pz{������iz]��#pw3��F�ߠ0b�rqY���;�BGm�.Ol�l<���������c-�i5�)��^�3VTm�y��Z�B����ӽ](��ȼ87Al�M1-�ə+��><a�º�0o��k���mZoL,P§4�TX�G���\�4�?V�ޒ����_fNɷ qz+j ��C�'����!�JmR�$�O�uI#��i���W���p�Џ�OHw\J��%�|̑�T��+z6Z]�Fy=���(0��O;8��C�Lm�V�{��3BU���2'�4K���~�4oL�d�;
� ���z�;�x�g���V��j��0=�P�jV������ɾ�]�E !�R�xs~[X`��8��AR���?�#���[W޾ҁ>�����1!�`֋8v�:hb���?\P��~r��Vw��j�[�go<��j�\a�e�Ȥ�?�/r�v�7e\�5�֎����r��Pw�R�h���fp �M����T%J|��8�ǩ*x���LJ<�F+t�`��s��$�fZ�.�E{+���4�����������ّ#�~�(󣛳���hP��&�i���G�b�5О�W��u�*�9�ע��,��:����M_�HY\C�@��FW�����Ɵ�fxr
�1���E������
�'�w�ӈf�{u�{�\��Dw��R��%xY��W'Aa���?��r�읉�Yd��^,�C����)aɺiP���NZ$p�s���-d�U�ȧ�o�P����Y%dZ�	o�7�B%<�C-W��8��Hq�����u~�6�>�?�ZM��&�]հ�����U�k�u�? ���s>��l�@���t��M�//!���z�HS��/�?zn=�����	�x3���in�b&�~�E"\c�k]���iJq�/t�;�j��k[f�~�U�'������M 9���M�{P� }RF7��b�Lp����JP�|d�C	����OIku�E{��TG��S*쳔��Lr��x�ʏsKb�{ ���݆��f�O���:�(qo���Y�1�9̓���zv�9D�`u��p�����p����a*���p�r^_��ב�_���j��Cޯ�:�/b�2�f^����ռ���p�1��ؤ����t���'8k�h��D����
 �� 9�$���� �'�ɩ
y7���:ĵ�c�gn-�O�.�X���|������r)z+P&�8��3`8����juŠo�.����E���ՠd�O��\~+gݪ&��y�- ��c,$e.:�ȁ��i���]v�+s�t������F�%J�6������%�\��'�bO��<��M�:�����b�n$���չ�;K��'��7{0�����ij ����"�5��VB, �l8m��,a��B����Ac;s�f��F�B���gs>w"����I�Si��N]�-nJ	�l�iK^�o��Qg�d��qH�ˌz&i�1��_6dN{=<O'��C�V�ů��k���U�]�l&�^qz�<�_�].�:�+ ��H'~���#��|�n��I��%�x��0���7�����z���Y� �8�8�F l�~��
��o��s�{ba˽����2�򴲁G!m�[���x�E�4j�ҶBO!�B�
��	��l+���$��7����]5t��r螔���	�#��Mo���CZ%C�^'h���*�Q�	9�b��+*P(���Yxx(��	�>d:O�IZ�!��u���@���8���ޛ�DT�CY�M]���O�dQR�aE�9D��]}G�v<b�ɿ��&j�svE���,�p/;��Pү}��O�?W�~`�d6�T�����)cyU_����V/^���o�I��[��6fL)����Ki��#fhO��u΢OW*��M�$`��Zf$� ��`�+x��ɇ�p�R����3NqߑHl@���G�g�޲?!��پ)^�?��,���Sz���P2!�W�Gaj. �k��@,��!�6m8��|M�'�\O������;���-z*��^��Y�u���Ό�_���Y���$3����|�\6~�G��~*-t&X�|����٪6����|��9Ũ�6�DgYu�YeG���OM(Ɲ��̾��G7��NQa\Bb��q�W"����R�^�󹳽�)��9z��s�rXO#I0%���\M�pte�e�ġ;n��?�����ߵ�KC�`�VTK����=��O�� �k:N�P�K"���w�?{�"�Q�C"t�CV�����?��S;���9�.��n�M���?������ "���~����p=ҜW���cx�c�-+���2Cy��ņ�%-��Q���q��3
�;Ф�ֻ� 8�Z� P�}�>m�8�f.��L{�����7Ъĝ8�)�6�ڛ�z��M/��a�B)�s��q�~�H�B�i�~����Ƈ��9�"�?핫g�����/�*�8�_�p�MWv�d�B�jy���B����GQ��	q�R��ߴg�k��zp ��Y�n����܉�"�T�ϯ�U�Jj�0D#	��Ϳ���->�>��˫	�cF�@��*(�ԇ�s�7I�R�`'ͪ�}��f���%8P��!NI��P9�oܡ:�oB��'�t��T;���V�\���C,p15)���r�W���p�[��%��ga�S(�k�c	���=�2��2Ӱ����m@mkmәXʧ�s�M�o�rn��C�LK`by/��u�{	��I�~΢6��tfw�=C��7��M�Kb/����τ�\*W���(~�V�_�6�wmvن�, ;�Q�p�7�� ���Ww����KzY���b�0�\,��Kq�Jo(}���V!��*��x')�P��qD'��</��Y�Č���2О���{fe��Y��!U[*��t�N��}EO��E�1�]Y^�Oa�C�� ��E�@�@�x�х����ǈ����U���]�X�&���2�T�P+����,�|����_�*�l���\4bk�B���7�Э�N����)ԅ:��q�>��m"C����Lq?,�����ГSo���sD<��VE�+0�Q�mFUyH��|J�ڔ!�o���U1�)O��������/���Zi�>���O܈�x���F��}��1�Ǚi�@��M$�DK]:h8{��TBWNO�Lp�����ý}.'�8�8�9�{�p�;�4H���'FHf|t���dqXvR��=R��V-������Bv���r{0�-pX��ml�Gu����&�O��ኗ�<����E��̴>Zbh?�b��V���Z����͕�_@iyS�"��w���2��'B���^��Ce5Y���!X>��&,��g��u�ؾϼj�ٮ�7��rO�3�d ��'T)�?�j�
�i�'P��D��	�ƿ[,2!�"{,fa@�a��<bW����R|��FD�R`�E"iÃ�ɊBG��p�1+���J��e�m&�ͧT�fa�G)<�@�:9�3:q�ݸH�_�u���L]~o�tj�cmڧyl����φ쩺�
�?��c^�_x�ܕf1��S0j!-?g�Gl��{e�TR%g�`6�-g:g��G�`�+u�G��O~M�{=���Ӑ���YqBR�&��5�D,�C���-{�≯{ֳ}�f�lD��pΠ��X�c=�n� �ۄ�q&���� J�G�Rڰ��)gߓD�,m�B�֎�Y���zC,�O2�$�p	�c�U̗6���X�y� �,�?��Q�I�e��z�Yݸ��siő>j��Őo�A@@�閡�YK8�5���<J�D�r�M���sz:�������.�Fg+����[R�@UW�ոM��_�P��tB�Zl(��H�Z�@pf��0�'�6Ào�!��^:����Avح���0jx��R���Uo_�z��&�m��]�y�O,w�։V����>�P�h���bG�M�wL�O��tdܾv[s�o�D�3'E�M�w�
~�HaYYi��m��C)̌x�{������Q8yE�mu)m@��3�� M��#���be��ل6G��e�y��(���r&T���L6����J���h�2��"�1��E.�����r�Q㉈���
��1��v�`Mii�����.��`�
	�"�48ʖ{$�>�7�Y�L�D���O.l����p?A�.��
��Ҋ����ŘR�2~�*t>�S��;Y�����DC� ������Y�lR����V9����3�3\�7��]���
KOj�E+��M��F�bvȣ�dҽh�X��
0���O'��P�e�^̱}��^��Ѵ*N�m�����FZ�S�`Δ%9�ݾ��ʇ$��i�p���}ǉ:S��8�`�-��>��^��0�Ç��W������F8UkL�T,�=R�����+mi��q��};@3�	K����P�[%��ϝ=����C�#��]qIg��#�v�/��pt>Hϣ&u��vD3r��&u��Dqz5���Q}h7cF���\g� :hpa�a��r�L	2��D�%����5�~z`�_�&V�)� �8Q��*�`<	ai�C����Wӣ��4V�w<뮤d�f��@��_g�x�MּX~�̴�/@�?laV�d�\M�-,�/���r��΍�ƷY��
_�<\�/�MK�]� �֧�q'�3J�ӱU�}��y�-~5gm�K�ZC/��Lq�ݦ���aaYW��d(K$H�v���.�$��7Q����A�nu|���͟m����xe�1D��4�G��=�)�s7]c��E  ���}������M�� �Ϸ�(��(Q�Ɵ:���p�/Փ꤃�sC% �����l̡������nW�]����O�G0���=����Kx��@������`�N��*iKњ��߉�r}��1t^���'ۇSטY`e�Q�LSl�)����(��S�l���e��q�OX���`���s�0�*�q��msr��s�%��-Tp�NR�e�)���4^ʗ.��¿��I[�ܲ�D|+��?	���z��uo����K�5o���h
3{^uM������&�9��%J�J�$�k<��~�|}ښ`G��/7���u�,l�2�`͸�C���:Q�3�@S�Q���t���؀��-p��A��3�ȼW�T�"�ǸRQ��/x��
�����W���_֠-p��%1!�U4I0�`��2����y��ﱵ�}U�-�^'9`�%2WZh��֜gƨ�m�e�#ʯs�U5oCزpة0K�7��Է�3
�y�g˘��BE��/A Q�C����� ��!a��k��n#9�{}��Ups;����	���W%��]\BҪ�#���qbb/��s��O���``���q	�O(-�;����7�7� �����(���WM�Rc��=��/ӉMX����0��k�M��=�{lA��JZ��#�L0�i$m$�zR��k5��՘��gA��"�U���1��Qm"�]��/a�c�a��tEF�1 �A��{e��N��&���>#d{i�<�Y#�uu$�"Ǹ������WN� �Y�R�U�2�o%�B<�W�i�ؒ�{�jh�\l@@�?~+��s�2��,���F���W^���7����ۿ�ߪ��jX���`'@���v�KhH����@
�.��삆��x2]������8�Y��4�6����C?�g����7dsC�PҜ�h��R{=V�թ�:��w��ǩ���e����"�?7��c��8@+�2�^��%�ͼ�a\jw��kI�8�R�#e��<�$.jo\�j��aʠ
�ør��Ej��!���slj�jċ8q�~��f@"๔���/�NT��� ���u�峺���O�nZS���ݗ��Ns�������|�U��9�w�A6����S*�N�yɎ���-m6�$�o���;%���/�ܙ0�"a���_�*g^i�]�r��p���%�x(�pH��Av�E4D���Y�(��~K�DQe�_-�n�aUݭ�
��Җ��@��&�DQ%Cɱ�h�6�C?�]�X�
}ZG���^�Ox�\ �|�7%I�	��<mT�g@�d�� �8$BS�!�<nh�8ܧ��rܜz�'��r �ƾ�V�t�b��s�WVq��G9�5��F���S�t-�&�*Wt[^������c��P)#�ߠ����&9�C@@8AUltG���䵠���VW��vZE���{c�a籮߸��=2�wv�~j�����Ԣ�0[�0�An{@-�\��(3[k�eI��ϐ�K�].ܹ�g~��W���}���'P�R�ytZ�O"}���#S��7�b��vk�m+����:_�Sjk&
�Qp��~����r�8އ��)g@��>a,!����D�㹼_�B)M�S�^,��^"�D�w����Io����^��5O����\������K�M/j�U�m�I�0���\�c�؁��l7��Օ�-6�����.�`�Y	H/
*M<�}稔�j5~HӬ�B�x6q[�5P�.ӱ'����3��i>-ޠ{g����lDu;�f��o��GoTV�u'{"q�Y	8�0!4	z3�r%s�6\(|�=� �t�\��6ӛ�d�)s���������������`L��Ǉ{2�]r��|��&�WSqVn�Q��=�����+n{����i̧G�ZZ%ʍ��Q�V/X�2��IGJ���>jF��5;I��+D�~f�T�쌩�*�p�D��fH��N@�T9���1�ND+��Kh�O7�/ٺ;B�?(R{<�O��PT�A05�57�l��C��0�����Φ+.�&O]c�JO�QS��TH8���ax��3Nj&����ɨ�͏����ψ���c`��Ďm��P4�+��9$��-%�W@)���3�{�T�B�\l��x8���ǙZ�L�z���F�,��'���t/�K�,��p�gNsw�Vc�G�]��a~�x׮,�;g��᠉C�1�/_j,	�QB{t����:��Hs)(���m��s�nٔ�7	Aq�-�mʏ��II쐹���EdF�#)e
��dK� X��1d'��G�U����ޘ���P��h��� ��g��)%�X����j��&�;f�I�ߙb:����+��ko�`��N����a��	4@�=v!Э����&�L��ջY���8��/��"��I���t��̯C�T����љ
�+}'��RÛ��~�\����>A�pZ|��)�B�[V;Ss�l_%7�i��8�q�x�E�RE���`�-���`m39�J!�k����1A��0�`f�,��_��J^���q��Xh�O��}=��z���;���itX��C(��Q�bH�~�q)����(�B�as��&x^��,"�̖�v�]a�̽wmRL��\ 뫵����[����U�QJ����=BP@����F�V�Y�9��,;[��ĥ��J�1����o�ӆXMab��H*F�B�N������@�πs�Ā-z����	�{\)�˵���Xڒy-�b��M��xT$].��ܺ y�.��RQ�_��Y��n��`���Ԟ���=�1刌�0�����K�cO@����8>��y�U���.!�$q�K�9Cr��~'"��<O�YD�@���.'a�u�[��j��)���������@&zVIX��y���*�:|���o�n����_q2�r�������X�9JR�X,:�m��DAHm�F��H�7�h9�Vn��L���cC��"e�=(z�a����kߕ�"�ɉdɂ��A8��Jq\���b�Hx����v��H��V�*!�=F��<N�$Ai�ق?��٥X��B�� 4�(q�M�9i*�X����FՂh�_�N�E�����aŰ���xc�:oU�~�.��Pk�����m��9�4�}!)Cm�����~k�c�c�pIYs|��᭒=29�1Ү�:��$.q�S@��*�E.!l��1X�2O���>���~�|�wy�����}��֫}�D�կ1T`D	�	eJO�d�& e���R�,�[���z"ıu����D�*�K�TndJ�6�9�6�l�O0�w����h<���0�h'�mH�1�=�D%�7
�{�����j��]Ï�87T���,qhBO�:3(k���_m��〪�=�-^��Hs��4՜������r�H�ST7�����G�b�)��h�u��/�7ψ����z?���1�1J���*��R5���)p�ڿ=�s	6���,�ı�������[�C[����7H�����;'%r��:���C]	R��+ �*��GL�#�8�7f��J�M��P!Pp d��B�#1���K�����pK$RW�*sj�*wv[����,u+VoT��[�FU��V)��R�i6"��s�������9����An�B�����>j���#�Yefey �u����Q1��T���ۑ��h�hF�����4�:�N;lcH��d�#/Ԩ��6��\.������{�����"Ggf�*��Ĉ��^�c�*�
<1A��6���;E�^���Վ��'�FԆi��E�+���3Uapg�bTGY��q��f{>�����zي(SUѯT]��o����T��ōh_}0ƽUw^ܼ����jȫWjTi0��j@K`�:$S&�ʁ�K��o�[�!L2g=����t/�m7��8�3n���3J9��ٓ�o��sL8y��C�=
��#�9F8C�YU�����{�H�����T�3�a���a,B���ыXH�o⣦��#E�^�z�	��BNjaA[��c^rH2��� Xp��\�H^ضc���4G��!��E��Ⴋ"-���T�6�Sj\�I��v�+k&���({�.;2B`����]ò��b�L}԰%� R�$�2R�Gos�Թz����?3�3BآvR=K�;q<
����?�������,"����!�G�@�;S_���X�G���eed��+��]߰o��&�*e���^.�WK��>��מ�A[!K(�z�D��p�����tI������#_��Z �5X�(6U۬F�"� h���%���Pi��1b��,�ZASL`�ҡ٥��Uj:8��0�,��N�We�Y4'Bmk,�N�с��啕�CEN��l� ���l�Hj\��-�)_��k���H�H'�9�*3D٣Z�^0�[v)`O��zR�u�,�D߯��|v����6�ؼ���%q=K�;;=F�>�Ԯ�?����}cC�uH�~�fV#���>���D3\���F��-X�w*7ݢ� �^�D�b������� 5$im���X&Z'���m�yu|7yt�����"��
\�P
������@
�$�W��;yM�3𽙔G�ˠ���� UN�����ɘ����R�<�!�7�)I1m��'Puz��J ��.�u7�;o]�Aw�(���^.����)�K��F}=�S��Q�|�ǿZ���K?Ny��؋Z�u5�����T�آ_!�/=�×Ek%�6ۙ�UA�P79&M���iHDz���M|J�W$V��>�C�B��ϳbj�~h����z��\���V���
�d�z��� �kya�����]��+G&]Bl��w(��	�˴:��r	��(��eFf�(���	f����*��V�^�~Q���yT��}�Q֧�yn`�1�*�@��2 HsMG&���|�o$N�ͥ�~��q�܍űs`���a�����MJ鰋��D�Ơ
�?o�Xx���a�5@���_�$��Ctw;�s�G9W�U|i�Ɂ���,O�| 7o�^~�MogZ��������M)Pn�����L+R��4��%�q�`�aȹ�=���f�LY��).n��W�Vv3�"hfNG��%��a:����p�Y}8���Q��wMIn���On��/	 ����J�ل���p?4��T���۞K5�,}^	X��%P��>u�P�=,gB��,�8&�A����'P��$�MM��r�Z�ڔ�f��q�U	���Ht2b�+�d��B��r�@��N*֊p�w�����!"��޿7�v+kP�7�n�kw�yF
���{<�:Hh�AgI��ͳ��U�=�W(kl}�5	<��S6�8r8�Z ����v��6~�ˠ8�ٮ�@�A�g�C�/�����sٍ2$^0��L�0,��[��j�J	a�O89���l!Q&�<$�:>A�3�px�g�\�a������������~Oˣ����gԣX!6�/8�]4��<d5�k'��O�4x��Ļ)�At��B�l{Y��ζ�#��Pyb�<�,k�/�M'X��q3d��h�}Sk�=D9g�Q�g�8����K�E�`~u�	4*@� Rv4A;z�L�Y�N���G�z�k6�(t��CH!s�da%}jS|r�_ղ�c4�(`{���!�M�`8���AqlE�{��N�!fq?�����SJ	�����Rg&�|A����/V�DK\Akl���綗���Y��򕍏*�·J괇�l6Ε�B�ۗ`��]֯��&y�E���L�4�H�[l�"��<G#	��E8��w�g���5�HM3|~�L�p�F���/�QC~��/��Xs��v��2�{;��¤�Ù���^d�Ӏm�L3�H	��}Ǭ?[_��J_�P�c�t�\������Ȗ���A�~f��r�?%ڐ��VL&�z�I%�h���!x�Z���s�?!w���C��	��W���5#:��)��ɫ�\�*EU�i�Lr���h�~
7��9���RϻK�4� I����3q�<Cf{M%���U���H��`#7�= H��1�n]���}c����R����CA����M:x�����\�������뎒ff��f-H�u�mW�[��}�(D?�/$㳉	(�x�����?��e���hWFR�$s��OT�>dt
d7�)�t�*/����d��E�&p��7��*��G�jŠY�u���%�����<8ʒp�ҘL�#<�%_5� 9���V
�+`נ�њы�h��A�?`��L�?�ҷ��N�o�TW��������B�O��I�>�$�Z-�?�VL-rI�$�'E&�;���*cS��]��3G�
�`9\2�A��9)�1CI_v�i��;��i�3&P�����AQ�1�_�-'����`�!�]�,�1,#, �}`{��s۵��uc0�ߟ������S\f�I-�n7j�_ke����7q/5��9��*k:�^��[��� ���4��VH��$�ƀ���Y�i�Z�V�)�QO �%�G:���b>ɩTH{;�Ϣ+�ŵ�T�	�-���6ק�igOG�0�Z�Z!���U�s����P�1/�^���\Q���	�x#v���)�K��^���*\���!�&�V>�)@ᴣja�%dc�����o�A ?�1�ބ�c&�u�W����SIh:��pf��̍���/`лΥb��@��H�T��Ɂ=Q�X�Qr���q2�s�=��/Þ��cJ��'���\�;�^�v]8A���")�R�7Ⳡ�D�]����j�蒑��r���|9��������r¯i,`�U@�A��T�6ע�5�v���Ot�I�-��s���E�׶�Zz?�0�n ,��}>����	7�M�}I�g�nX�O�H��O�S��Q��|hQ� >w���Sx�	"�3��#�[bDt�d�8S���S�����5�2�d��m�B�vto^��c���4=�ʎ[� ��$[��Q0��ˀ�>��������N:D`ƒ۽r|,�����<����fe�t��ۓ�
���V�?�LŜ���J�O�1]V�h�c�z(l4=�_Q֌��ߎɟ�������pu%�
���I~��Uhmy�Nbi�AQ � 9�.��Qޗ@�
�Z�78�w�� �����zw�9V��VY�˳��8A�nd�L���\;	���/	,$��k=M��s�����
���Q�m�r>� ��Y�4yЕ�j�r�����x/��WQ�v�{/��{`:�/��,���8��rZ_o�������o,���;$�b�	C��4ׄm�s�D�[НVkb���a&�Q�ܜBM��R��x�_�g�9�LT�Hd����CjS,�rf��r��U�Tk��6E�-����������7�,ZL���մ��f}
Ɂ�)cL���#��-�z�Xm�O*�Nd�����a�o�s<���9%9>�o�,{a���E�UQe�	�qC:���1���S+#1�¡]�o���BQ�J�޵�stx��O�Y�UP�a�KR���W�r13@��i�^�-��.	
�����^�/�z�LV�x��S��%��Sfw����fJ�����ˉ��n�C:��4
B�|GD����_85AvB6~>����?s�n9gEF���������Xq�c�p[���qŽXEI�W��p��SC���Pz��������1*s�^o�����z����A��l�� �n�Fd	���σ�.�D�w��^8�D�.VĊ@I�n��a��U"lY����ӎ���ڹO	��;����1�B�=���L/����`"�'�<���Z�7��e�3�jY�����ςa�R���z�y�
T�M�O�st&@
�9螄�x}AW�zw5gȿUy�_GР*I뭼+�����<l_p�@�nyn�P"����)�3gɇ4L���!ƴ�j$��ς:�玕p�պ�ncf�������{�ֶ�ۣ�˥a��߁yoG��֡L�$��Hgٻ�x,���H��RH�:�q���2�����M$���Bۚ{���P�y�{�G�>�N�;�:k*��� f��>$)e���r��ǝ�-a�5�&B[�<�������]��5�sC��:!�U�!���lFm���9���&Y�[��|L%V!���IF_��
s�B����rXP�5������q��<L��Y�l�W�z���Ct���������X��GPs1�������{t�W�{�X��8U����K��w��X�dM���8�eyDL���#I��NVC	��yo��E;�|�?^Rx;	�$�D�n3�y�n�\f�BeM�6A�R��Vp��vy;_痢�]bĠ���M#��*�m��+��^(E�^��������:k��!Ք�i�cZct
�a�H�� iA�N�ժ	T�C�*V��ƀ���leL�z�C�o*n QR�E���:�%��|�,�CԂ�5�Tu�H�B.î6T8�N��ǂ�HXz��l�žk`��=R��2�\w:o���:�6�&մ�f�f�j�Zi��I���0}�A�7jQ�q��(Iydh�h�K�f�`^�����r��۬0W��q MJR������y"�]��`���֝j�����OH@���<�n���ީD�(V)�T#�Z�"6�2Ґ���J����Ҏ��(k�a5�.��tp1~q�>^��QĔm���X8Nh�%8T�Bu���l�BzS�Z�x5s�� �cV��X%��g^/�UN��	���-���1����|h^3�J�'�O���~���a�1�y�x>O�0ȶ��rʺ�U����z�I��m}xJ��p�����Nd�եJ�ut�?f��2˾�(̅\�~��1fO�FN7%���'��&�a��{�����f�֜cvvn[b�������{�b�T�>���[,	aP�!�)��!�{�69����-�qF�P�*gT|<
�8z�����
Sj�*��7I��y1�w�S�~��&=�J�T��3�<�/��س{ž �9��B8`�'�z�c�yἚe>_�[��h��RN�2�Mà��HgC�ST�[á��Y��:Һ����k0�_�m�S(M'5tx�8�U��"v)���4�"�Ƽ��<g(Ӌ2���Mf�D��F�#����-��.כ�xM9`BJޤ��7:UV�8���.@)+:�|W='EfLj����2XLyC���aܬE��?�צ}��V��`�խ�V�uz/lؚ��ӎ�IZj�4/�n����C]$�s�����V!!�-b��\'4�QZ�D��
3.A���t!\���ù��m�b��Q�S�����Y�
���-�?�"���w_�"�x���� �&���Z�#��@N��A��u�~Oa�;�D~AT
�u$�y�)*pÏ|����&Ŧ�(wx�@c�N���u4�m"h%�79P Yhz�}*L#^X���9OŰ%܇	�0h���Q{IK�s�3��'�״����͊F�I�����P��^��:�'۳9���4wL,R�0aT�(����P`��)ٞ�7�"L��
 ��7��/���'5E� ����?C�S ��N,��I,x/c�r�m.iSY@��87�0__kl!�^�H[�,�!:�c��+f��լ,Ŵ���$ ��?��S��6���,XbD��sC`I������I8��e.�~	�ކ8�@-Tih�9yЌ��TW\o������V��a͠�խ�oES�#�G|
�?�:�Nk�M�I���Q�Ά�$��"
W����ж?��#(�	�=V�l�?��4^w`+N��;uF�p�V�o��[�v�2ｿx�����1M _w@��L��{�������Ooh.�/7�	