  --Example instantiation for system 'processador'
  processador_inst : processador
    port map(
      DEN_from_the_lcd_sync_generator => DEN_from_the_lcd_sync_generator,
      HD_from_the_lcd_sync_generator => HD_from_the_lcd_sync_generator,
      RGB_OUT_from_the_lcd_sync_generator => RGB_OUT_from_the_lcd_sync_generator,
      VD_from_the_lcd_sync_generator => VD_from_the_lcd_sync_generator,
      bidir_port_to_and_from_the_lcd_i2c_sdat => bidir_port_to_and_from_the_lcd_i2c_sdat,
      counter_from_the_fft_pipeline_0 => counter_from_the_fft_pipeline_0,
      ena_10_from_the_tse_mac => ena_10_from_the_tse_mac,
      eth_mode_from_the_tse_mac => eth_mode_from_the_tse_mac,
      gm_tx_d_from_the_tse_mac => gm_tx_d_from_the_tse_mac,
      gm_tx_en_from_the_tse_mac => gm_tx_en_from_the_tse_mac,
      gm_tx_err_from_the_tse_mac => gm_tx_err_from_the_tse_mac,
      local_init_done_from_the_sdram => local_init_done_from_the_sdram,
      local_refresh_ack_from_the_sdram => local_refresh_ack_from_the_sdram,
      local_wdata_req_from_the_sdram => local_wdata_req_from_the_sdram,
      m_tx_d_from_the_tse_mac => m_tx_d_from_the_tse_mac,
      m_tx_en_from_the_tse_mac => m_tx_en_from_the_tse_mac,
      m_tx_err_from_the_tse_mac => m_tx_err_from_the_tse_mac,
      mdc_from_the_tse_mac => mdc_from_the_tse_mac,
      mdio_oen_from_the_tse_mac => mdio_oen_from_the_tse_mac,
      mdio_out_from_the_tse_mac => mdio_out_from_the_tse_mac,
      mem_addr_from_the_sdram => mem_addr_from_the_sdram,
      mem_ba_from_the_sdram => mem_ba_from_the_sdram,
      mem_cas_n_from_the_sdram => mem_cas_n_from_the_sdram,
      mem_cke_from_the_sdram => mem_cke_from_the_sdram,
      mem_clk_n_to_and_from_the_sdram => mem_clk_n_to_and_from_the_sdram,
      mem_clk_to_and_from_the_sdram => mem_clk_to_and_from_the_sdram,
      mem_cs_n_from_the_sdram => mem_cs_n_from_the_sdram,
      mem_dm_from_the_sdram => mem_dm_from_the_sdram,
      mem_dq_to_and_from_the_sdram => mem_dq_to_and_from_the_sdram,
      mem_dqs_to_and_from_the_sdram => mem_dqs_to_and_from_the_sdram,
      mem_ras_n_from_the_sdram => mem_ras_n_from_the_sdram,
      mem_we_n_from_the_sdram => mem_we_n_from_the_sdram,
      out_port_from_the_lcd_i2c_en => out_port_from_the_lcd_i2c_en,
      out_port_from_the_lcd_i2c_scl => out_port_from_the_lcd_i2c_scl,
      reset_phy_clk_n_from_the_sdram => reset_phy_clk_n_from_the_sdram,
      sdram_aux_full_rate_clk_out => sdram_aux_full_rate_clk_out,
      sdram_aux_half_rate_clk_out => sdram_aux_half_rate_clk_out,
      sdram_phy_clk_out => sdram_phy_clk_out,
      tx_out_from_the_fft_pipeline_0 => tx_out_from_the_fft_pipeline_0,
      clk100MHz => clk100MHz,
      clk50Mhz => clk50Mhz,
      global_reset_n_to_the_sdram => global_reset_n_to_the_sdram,
      gm_rx_d_to_the_tse_mac => gm_rx_d_to_the_tse_mac,
      gm_rx_dv_to_the_tse_mac => gm_rx_dv_to_the_tse_mac,
      gm_rx_err_to_the_tse_mac => gm_rx_err_to_the_tse_mac,
      m_rx_col_to_the_tse_mac => m_rx_col_to_the_tse_mac,
      m_rx_crs_to_the_tse_mac => m_rx_crs_to_the_tse_mac,
      m_rx_d_to_the_tse_mac => m_rx_d_to_the_tse_mac,
      m_rx_en_to_the_tse_mac => m_rx_en_to_the_tse_mac,
      m_rx_err_to_the_tse_mac => m_rx_err_to_the_tse_mac,
      mdio_in_to_the_tse_mac => mdio_in_to_the_tse_mac,
      reset_n => reset_n,
      rx_clk_to_the_tse_mac => rx_clk_to_the_tse_mac,
      rx_in_to_the_fft_pipeline_0 => rx_in_to_the_fft_pipeline_0,
      set_1000_to_the_tse_mac => set_1000_to_the_tse_mac,
      set_10_to_the_tse_mac => set_10_to_the_tse_mac,
      tx_clk_to_the_tse_mac => tx_clk_to_the_tse_mac
    );


