--megafunction wizard: %Altera SOPC Builder%
--GENERATION: STANDARD
--VERSION: WM1.0


--Legal Notice: (C)2012 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpuNios_jtag_debug_module_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpuNios_data_master_debugaccess : IN STD_LOGIC;
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpuNios_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_instruction_master_read : IN STD_LOGIC;
                 signal cpuNios_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpuNios_jtag_debug_module_resetrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_granted_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                 signal cpuNios_instruction_master_granted_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                 signal cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                 signal cpuNios_instruction_master_read_data_valid_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                 signal cpuNios_instruction_master_requests_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                 signal cpuNios_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal cpuNios_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                 signal cpuNios_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpuNios_jtag_debug_module_chipselect : OUT STD_LOGIC;
                 signal cpuNios_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                 signal cpuNios_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpuNios_jtag_debug_module_reset_n : OUT STD_LOGIC;
                 signal cpuNios_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                 signal cpuNios_jtag_debug_module_write : OUT STD_LOGIC;
                 signal cpuNios_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpuNios_jtag_debug_module_end_xfer : OUT STD_LOGIC
              );
end entity cpuNios_jtag_debug_module_arbitrator;


architecture europa of cpuNios_jtag_debug_module_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal cpuNios_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_instruction_master_continuerequest :  STD_LOGIC;
                signal cpuNios_instruction_master_saved_grant_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_allgrants :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_allow_new_arb_cycle :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_any_continuerequest :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpuNios_jtag_debug_module_arb_counter_enable :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_arb_share_counter :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_arb_share_counter_next_value :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_arb_share_set_values :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpuNios_jtag_debug_module_arbitration_holdoff_internal :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_beginbursttransfer_internal :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_begins_xfer :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpuNios_jtag_debug_module_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpuNios_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_firsttransfer :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpuNios_jtag_debug_module_in_a_read_cycle :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_in_a_write_cycle :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpuNios_jtag_debug_module_non_bursting_master_requests :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_reg_firsttransfer :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpuNios_jtag_debug_module_slavearbiterlockenable :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_slavearbiterlockenable2 :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_unreg_firsttransfer :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_waits_for_read :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal internal_cpuNios_instruction_master_granted_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal internal_cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal internal_cpuNios_instruction_master_requests_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_cpuNios_data_master_granted_slave_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_cpuNios_instruction_master_granted_slave_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal shifted_address_to_cpuNios_jtag_debug_module_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal shifted_address_to_cpuNios_jtag_debug_module_from_cpuNios_instruction_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_cpuNios_jtag_debug_module_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cpuNios_jtag_debug_module_end_xfer;
    end if;

  end process;

  cpuNios_jtag_debug_module_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module OR internal_cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module));
  --assign cpuNios_jtag_debug_module_readdata_from_sa = cpuNios_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpuNios_jtag_debug_module_readdata_from_sa <= cpuNios_jtag_debug_module_readdata;
  internal_cpuNios_data_master_requests_cpuNios_jtag_debug_module <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("100000000000011100000000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --cpuNios_jtag_debug_module_arb_share_counter set values, which is an e_mux
  cpuNios_jtag_debug_module_arb_share_set_values <= std_logic'('1');
  --cpuNios_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  cpuNios_jtag_debug_module_non_bursting_master_requests <= ((internal_cpuNios_data_master_requests_cpuNios_jtag_debug_module OR internal_cpuNios_instruction_master_requests_cpuNios_jtag_debug_module) OR internal_cpuNios_data_master_requests_cpuNios_jtag_debug_module) OR internal_cpuNios_instruction_master_requests_cpuNios_jtag_debug_module;
  --cpuNios_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  cpuNios_jtag_debug_module_any_bursting_master_saved_grant <= std_logic'('0');
  --cpuNios_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  cpuNios_jtag_debug_module_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpuNios_jtag_debug_module_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_jtag_debug_module_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(cpuNios_jtag_debug_module_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_jtag_debug_module_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --cpuNios_jtag_debug_module_allgrants all slave grants, which is an e_mux
  cpuNios_jtag_debug_module_allgrants <= (((or_reduce(cpuNios_jtag_debug_module_grant_vector)) OR (or_reduce(cpuNios_jtag_debug_module_grant_vector))) OR (or_reduce(cpuNios_jtag_debug_module_grant_vector))) OR (or_reduce(cpuNios_jtag_debug_module_grant_vector));
  --cpuNios_jtag_debug_module_end_xfer assignment, which is an e_assign
  cpuNios_jtag_debug_module_end_xfer <= NOT ((cpuNios_jtag_debug_module_waits_for_read OR cpuNios_jtag_debug_module_waits_for_write));
  --end_xfer_arb_share_counter_term_cpuNios_jtag_debug_module arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cpuNios_jtag_debug_module <= cpuNios_jtag_debug_module_end_xfer AND (((NOT cpuNios_jtag_debug_module_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cpuNios_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  cpuNios_jtag_debug_module_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cpuNios_jtag_debug_module AND cpuNios_jtag_debug_module_allgrants)) OR ((end_xfer_arb_share_counter_term_cpuNios_jtag_debug_module AND NOT cpuNios_jtag_debug_module_non_bursting_master_requests));
  --cpuNios_jtag_debug_module_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpuNios_jtag_debug_module_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(cpuNios_jtag_debug_module_arb_counter_enable) = '1' then 
        cpuNios_jtag_debug_module_arb_share_counter <= cpuNios_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpuNios_jtag_debug_module_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(cpuNios_jtag_debug_module_master_qreq_vector) AND end_xfer_arb_share_counter_term_cpuNios_jtag_debug_module)) OR ((end_xfer_arb_share_counter_term_cpuNios_jtag_debug_module AND NOT cpuNios_jtag_debug_module_non_bursting_master_requests)))) = '1' then 
        cpuNios_jtag_debug_module_slavearbiterlockenable <= cpuNios_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master cpuNios/jtag_debug_module arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= cpuNios_jtag_debug_module_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --cpuNios_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cpuNios_jtag_debug_module_slavearbiterlockenable2 <= cpuNios_jtag_debug_module_arb_share_counter_next_value;
  --cpuNios/data_master cpuNios/jtag_debug_module arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= cpuNios_jtag_debug_module_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --cpuNios/instruction_master cpuNios/jtag_debug_module arbiterlock, which is an e_assign
  cpuNios_instruction_master_arbiterlock <= cpuNios_jtag_debug_module_slavearbiterlockenable AND cpuNios_instruction_master_continuerequest;
  --cpuNios/instruction_master cpuNios/jtag_debug_module arbiterlock2, which is an e_assign
  cpuNios_instruction_master_arbiterlock2 <= cpuNios_jtag_debug_module_slavearbiterlockenable2 AND cpuNios_instruction_master_continuerequest;
  --cpuNios/instruction_master granted cpuNios/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpuNios_instruction_master_granted_slave_cpuNios_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpuNios_instruction_master_granted_slave_cpuNios_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpuNios_instruction_master_saved_grant_cpuNios_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpuNios_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_cpuNios_instruction_master_requests_cpuNios_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpuNios_instruction_master_granted_slave_cpuNios_jtag_debug_module))))));
    end if;

  end process;

  --cpuNios_instruction_master_continuerequest continued request, which is an e_mux
  cpuNios_instruction_master_continuerequest <= last_cycle_cpuNios_instruction_master_granted_slave_cpuNios_jtag_debug_module AND internal_cpuNios_instruction_master_requests_cpuNios_jtag_debug_module;
  --cpuNios_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  cpuNios_jtag_debug_module_any_continuerequest <= cpuNios_instruction_master_continuerequest OR cpuNios_data_master_continuerequest;
  internal_cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module <= internal_cpuNios_data_master_requests_cpuNios_jtag_debug_module AND NOT (((((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write)) OR cpuNios_instruction_master_arbiterlock));
  --cpuNios_jtag_debug_module_writedata mux, which is an e_mux
  cpuNios_jtag_debug_module_writedata <= cpuNios_data_master_writedata;
  internal_cpuNios_instruction_master_requests_cpuNios_jtag_debug_module <= ((to_std_logic(((Std_Logic_Vector'(cpuNios_instruction_master_address_to_slave(26 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("100000000000011100000000000")))) AND (cpuNios_instruction_master_read))) AND cpuNios_instruction_master_read;
  --cpuNios/data_master granted cpuNios/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpuNios_data_master_granted_slave_cpuNios_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpuNios_data_master_granted_slave_cpuNios_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpuNios_data_master_saved_grant_cpuNios_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpuNios_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_cpuNios_data_master_requests_cpuNios_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpuNios_data_master_granted_slave_cpuNios_jtag_debug_module))))));
    end if;

  end process;

  --cpuNios_data_master_continuerequest continued request, which is an e_mux
  cpuNios_data_master_continuerequest <= last_cycle_cpuNios_data_master_granted_slave_cpuNios_jtag_debug_module AND internal_cpuNios_data_master_requests_cpuNios_jtag_debug_module;
  internal_cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module <= internal_cpuNios_instruction_master_requests_cpuNios_jtag_debug_module AND NOT (cpuNios_data_master_arbiterlock);
  --allow new arb cycle for cpuNios/jtag_debug_module, which is an e_assign
  cpuNios_jtag_debug_module_allow_new_arb_cycle <= NOT cpuNios_data_master_arbiterlock AND NOT cpuNios_instruction_master_arbiterlock;
  --cpuNios/instruction_master assignment into master qualified-requests vector for cpuNios/jtag_debug_module, which is an e_assign
  cpuNios_jtag_debug_module_master_qreq_vector(0) <= internal_cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module;
  --cpuNios/instruction_master grant cpuNios/jtag_debug_module, which is an e_assign
  internal_cpuNios_instruction_master_granted_cpuNios_jtag_debug_module <= cpuNios_jtag_debug_module_grant_vector(0);
  --cpuNios/instruction_master saved-grant cpuNios/jtag_debug_module, which is an e_assign
  cpuNios_instruction_master_saved_grant_cpuNios_jtag_debug_module <= cpuNios_jtag_debug_module_arb_winner(0) AND internal_cpuNios_instruction_master_requests_cpuNios_jtag_debug_module;
  --cpuNios/data_master assignment into master qualified-requests vector for cpuNios/jtag_debug_module, which is an e_assign
  cpuNios_jtag_debug_module_master_qreq_vector(1) <= internal_cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module;
  --cpuNios/data_master grant cpuNios/jtag_debug_module, which is an e_assign
  internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module <= cpuNios_jtag_debug_module_grant_vector(1);
  --cpuNios/data_master saved-grant cpuNios/jtag_debug_module, which is an e_assign
  cpuNios_data_master_saved_grant_cpuNios_jtag_debug_module <= cpuNios_jtag_debug_module_arb_winner(1) AND internal_cpuNios_data_master_requests_cpuNios_jtag_debug_module;
  --cpuNios/jtag_debug_module chosen-master double-vector, which is an e_assign
  cpuNios_jtag_debug_module_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((cpuNios_jtag_debug_module_master_qreq_vector & cpuNios_jtag_debug_module_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT cpuNios_jtag_debug_module_master_qreq_vector & NOT cpuNios_jtag_debug_module_master_qreq_vector))) + (std_logic_vector'("000") & (cpuNios_jtag_debug_module_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  cpuNios_jtag_debug_module_arb_winner <= A_WE_StdLogicVector((std_logic'(((cpuNios_jtag_debug_module_allow_new_arb_cycle AND or_reduce(cpuNios_jtag_debug_module_grant_vector)))) = '1'), cpuNios_jtag_debug_module_grant_vector, cpuNios_jtag_debug_module_saved_chosen_master_vector);
  --saved cpuNios_jtag_debug_module_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpuNios_jtag_debug_module_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(cpuNios_jtag_debug_module_allow_new_arb_cycle) = '1' then 
        cpuNios_jtag_debug_module_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(cpuNios_jtag_debug_module_grant_vector)) = '1'), cpuNios_jtag_debug_module_grant_vector, cpuNios_jtag_debug_module_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  cpuNios_jtag_debug_module_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((cpuNios_jtag_debug_module_chosen_master_double_vector(1) OR cpuNios_jtag_debug_module_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((cpuNios_jtag_debug_module_chosen_master_double_vector(0) OR cpuNios_jtag_debug_module_chosen_master_double_vector(2)))));
  --cpuNios/jtag_debug_module chosen master rotated left, which is an e_assign
  cpuNios_jtag_debug_module_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(cpuNios_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(cpuNios_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --cpuNios/jtag_debug_module's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpuNios_jtag_debug_module_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(cpuNios_jtag_debug_module_grant_vector)) = '1' then 
        cpuNios_jtag_debug_module_arb_addend <= A_WE_StdLogicVector((std_logic'(cpuNios_jtag_debug_module_end_xfer) = '1'), cpuNios_jtag_debug_module_chosen_master_rot_left, cpuNios_jtag_debug_module_grant_vector);
      end if;
    end if;

  end process;

  cpuNios_jtag_debug_module_begintransfer <= cpuNios_jtag_debug_module_begins_xfer;
  --cpuNios_jtag_debug_module_reset_n assignment, which is an e_assign
  cpuNios_jtag_debug_module_reset_n <= reset_n;
  --assign cpuNios_jtag_debug_module_resetrequest_from_sa = cpuNios_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpuNios_jtag_debug_module_resetrequest_from_sa <= cpuNios_jtag_debug_module_resetrequest;
  cpuNios_jtag_debug_module_chipselect <= internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module OR internal_cpuNios_instruction_master_granted_cpuNios_jtag_debug_module;
  --cpuNios_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  cpuNios_jtag_debug_module_firsttransfer <= A_WE_StdLogic((std_logic'(cpuNios_jtag_debug_module_begins_xfer) = '1'), cpuNios_jtag_debug_module_unreg_firsttransfer, cpuNios_jtag_debug_module_reg_firsttransfer);
  --cpuNios_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  cpuNios_jtag_debug_module_unreg_firsttransfer <= NOT ((cpuNios_jtag_debug_module_slavearbiterlockenable AND cpuNios_jtag_debug_module_any_continuerequest));
  --cpuNios_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpuNios_jtag_debug_module_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cpuNios_jtag_debug_module_begins_xfer) = '1' then 
        cpuNios_jtag_debug_module_reg_firsttransfer <= cpuNios_jtag_debug_module_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cpuNios_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cpuNios_jtag_debug_module_beginbursttransfer_internal <= cpuNios_jtag_debug_module_begins_xfer;
  --cpuNios_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  cpuNios_jtag_debug_module_arbitration_holdoff_internal <= cpuNios_jtag_debug_module_begins_xfer AND cpuNios_jtag_debug_module_firsttransfer;
  --cpuNios_jtag_debug_module_write assignment, which is an e_mux
  cpuNios_jtag_debug_module_write <= internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module AND cpuNios_data_master_write;
  shifted_address_to_cpuNios_jtag_debug_module_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --cpuNios_jtag_debug_module_address mux, which is an e_mux
  cpuNios_jtag_debug_module_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module)) = '1'), (A_SRL(shifted_address_to_cpuNios_jtag_debug_module_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_cpuNios_jtag_debug_module_from_cpuNios_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 9);
  shifted_address_to_cpuNios_jtag_debug_module_from_cpuNios_instruction_master <= cpuNios_instruction_master_address_to_slave;
  --d1_cpuNios_jtag_debug_module_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cpuNios_jtag_debug_module_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cpuNios_jtag_debug_module_end_xfer <= cpuNios_jtag_debug_module_end_xfer;
    end if;

  end process;

  --cpuNios_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  cpuNios_jtag_debug_module_waits_for_read <= cpuNios_jtag_debug_module_in_a_read_cycle AND cpuNios_jtag_debug_module_begins_xfer;
  --cpuNios_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  cpuNios_jtag_debug_module_in_a_read_cycle <= ((internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module AND cpuNios_data_master_read)) OR ((internal_cpuNios_instruction_master_granted_cpuNios_jtag_debug_module AND cpuNios_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cpuNios_jtag_debug_module_in_a_read_cycle;
  --cpuNios_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  cpuNios_jtag_debug_module_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_jtag_debug_module_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --cpuNios_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  cpuNios_jtag_debug_module_in_a_write_cycle <= internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cpuNios_jtag_debug_module_in_a_write_cycle;
  wait_for_cpuNios_jtag_debug_module_counter <= std_logic'('0');
  --cpuNios_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  cpuNios_jtag_debug_module_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpuNios_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --debugaccess mux, which is an e_mux
  cpuNios_jtag_debug_module_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_cpuNios_jtag_debug_module <= internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module <= internal_cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_cpuNios_jtag_debug_module <= internal_cpuNios_data_master_requests_cpuNios_jtag_debug_module;
  --vhdl renameroo for output signals
  cpuNios_instruction_master_granted_cpuNios_jtag_debug_module <= internal_cpuNios_instruction_master_granted_cpuNios_jtag_debug_module;
  --vhdl renameroo for output signals
  cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module <= internal_cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module;
  --vhdl renameroo for output signals
  cpuNios_instruction_master_requests_cpuNios_jtag_debug_module <= internal_cpuNios_instruction_master_requests_cpuNios_jtag_debug_module;
--synthesis translate_off
    --cpuNios/jtag_debug_module enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpuNios_data_master_granted_cpuNios_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpuNios_instruction_master_granted_cpuNios_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line, now);
          write(write_line, string'(": "));
          write(write_line, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line.all);
          deallocate (write_line);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line1 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_saved_grant_cpuNios_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpuNios_instruction_master_saved_grant_cpuNios_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line1, now);
          write(write_line1, string'(": "));
          write(write_line1, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line1.all);
          deallocate (write_line1);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_sgdma_csr_irq_from_sa_clock_crossing_cpuNios_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity lcd_sgdma_csr_irq_from_sa_clock_crossing_cpuNios_data_master_module;


architecture europa of lcd_sgdma_csr_irq_from_sa_clock_crossing_cpuNios_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cpuNios_data_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clk100MHz : IN STD_LOGIC;
                 signal clk100MHz_reset_n : IN STD_LOGIC;
                 signal cpuNios_data_master_address : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_granted_cpuNios_jtag_debug_module : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_descriptor_memory_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_lcd_i2c_en_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_lcd_i2c_scl_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_lcd_i2c_sdat_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_performance_counter_control_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_sgdma_rx_csr : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_sgdma_tx_csr : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_sysid_control_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_granted_tse_mac_control_port : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_lcd_i2c_en_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_performance_counter_control_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_sgdma_rx_csr : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_sgdma_tx_csr : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_sysid_control_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_tse_mac_control_port : IN STD_LOGIC;
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_cpuNios_jtag_debug_module : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_fft_pipeline_0_avalon_slave_0 : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_lcd_i2c_en_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_lcd_i2c_scl_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_lcd_i2c_sdat_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_performance_counter_control_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_sgdma_rx_csr : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_sgdma_tx_csr : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_tse_mac_control_port : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_cpuNios_jtag_debug_module : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_descriptor_memory_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_lcd_i2c_en_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_lcd_i2c_scl_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_lcd_i2c_sdat_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_performance_counter_control_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_sgdma_rx_csr : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_sgdma_tx_csr : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_sysid_control_slave : IN STD_LOGIC;
                 signal cpuNios_data_master_requests_tse_mac_control_port : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal d1_cpuNios_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_cpu_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                 signal d1_fft_pipeline_0_avalon_slave_0_end_xfer : IN STD_LOGIC;
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                 signal d1_lcd_i2c_en_s1_end_xfer : IN STD_LOGIC;
                 signal d1_lcd_i2c_scl_s1_end_xfer : IN STD_LOGIC;
                 signal d1_lcd_i2c_sdat_s1_end_xfer : IN STD_LOGIC;
                 signal d1_performance_counter_control_slave_end_xfer : IN STD_LOGIC;
                 signal d1_sgdma_rx_csr_end_xfer : IN STD_LOGIC;
                 signal d1_sgdma_tx_csr_end_xfer : IN STD_LOGIC;
                 signal d1_sys_clk_timer_s1_end_xfer : IN STD_LOGIC;
                 signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                 signal d1_tse_mac_control_port_end_xfer : IN STD_LOGIC;
                 signal descriptor_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal fft_pipeline_0_avalon_slave_0_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal lcd_i2c_en_s1_readdata_from_sa : IN STD_LOGIC;
                 signal lcd_i2c_scl_s1_readdata_from_sa : IN STD_LOGIC;
                 signal lcd_i2c_sdat_s1_readdata_from_sa : IN STD_LOGIC;
                 signal lcd_sgdma_csr_irq_from_sa : IN STD_LOGIC;
                 signal performance_counter_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                 signal registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_csr_irq_from_sa : IN STD_LOGIC;
                 signal sgdma_rx_csr_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_csr_irq_from_sa : IN STD_LOGIC;
                 signal sgdma_tx_csr_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sys_clk_timer_s1_irq_from_sa : IN STD_LOGIC;
                 signal sys_clk_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_control_port_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpuNios_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpuNios_data_master_waitrequest : OUT STD_LOGIC
              );
end entity cpuNios_data_master_arbitrator;


architecture europa of cpuNios_data_master_arbitrator is
component lcd_sgdma_csr_irq_from_sa_clock_crossing_cpuNios_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component lcd_sgdma_csr_irq_from_sa_clock_crossing_cpuNios_data_master_module;

                signal clk100MHz_lcd_sgdma_csr_irq_from_sa :  STD_LOGIC;
                signal cpuNios_data_master_run :  STD_LOGIC;
                signal internal_cpuNios_data_master_address_to_slave :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal internal_cpuNios_data_master_waitrequest :  STD_LOGIC;
                signal p1_registered_cpuNios_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal registered_cpuNios_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module OR NOT cpuNios_data_master_requests_cpuNios_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_granted_cpuNios_jtag_debug_module OR NOT cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module OR NOT cpuNios_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module OR NOT cpuNios_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 OR cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1) OR NOT cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 OR NOT cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 OR NOT cpuNios_data_master_read) OR ((cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 AND cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 OR NOT ((cpuNios_data_master_read OR cpuNios_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT cpu_ddr_clock_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_read OR cpuNios_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpuNios_data_master_qualified_request_descriptor_memory_s1 OR registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1) OR NOT cpuNios_data_master_requests_descriptor_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_granted_descriptor_memory_s1 OR NOT cpuNios_data_master_qualified_request_descriptor_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpuNios_data_master_qualified_request_descriptor_memory_s1 OR NOT cpuNios_data_master_read) OR ((registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1 AND cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_descriptor_memory_s1 OR NOT ((cpuNios_data_master_read OR cpuNios_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_read OR cpuNios_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 OR NOT cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 OR NOT ((cpuNios_data_master_read OR cpuNios_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_read OR cpuNios_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 OR NOT ((cpuNios_data_master_read OR cpuNios_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_read OR cpuNios_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")));
  --cascaded wait assignment, which is an e_assign
  cpuNios_data_master_run <= (r_0 AND r_1) AND r_2;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave OR NOT cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave OR NOT ((cpuNios_data_master_read OR cpuNios_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_read OR cpuNios_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave OR NOT ((cpuNios_data_master_read OR cpuNios_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_read OR cpuNios_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_qualified_request_lcd_i2c_en_s1 OR NOT cpuNios_data_master_requests_lcd_i2c_en_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_lcd_i2c_en_s1 OR NOT cpuNios_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_lcd_i2c_en_s1 OR NOT cpuNios_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 OR NOT cpuNios_data_master_requests_lcd_i2c_scl_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 OR NOT cpuNios_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 OR NOT cpuNios_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 OR NOT cpuNios_data_master_requests_lcd_i2c_sdat_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 OR NOT cpuNios_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 OR NOT cpuNios_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpuNios_data_master_qualified_request_performance_counter_control_slave OR registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave) OR NOT cpuNios_data_master_requests_performance_counter_control_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpuNios_data_master_qualified_request_performance_counter_control_slave OR NOT cpuNios_data_master_read) OR ((registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave AND cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_performance_counter_control_slave OR NOT ((cpuNios_data_master_read OR cpuNios_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_read OR cpuNios_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_qualified_request_sgdma_rx_csr OR NOT cpuNios_data_master_requests_sgdma_rx_csr))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_sgdma_rx_csr OR NOT cpuNios_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_sgdma_rx_csr OR NOT cpuNios_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_qualified_request_sgdma_tx_csr OR NOT cpuNios_data_master_requests_sgdma_tx_csr)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_sgdma_tx_csr OR NOT cpuNios_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_sgdma_tx_csr OR NOT cpuNios_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_qualified_request_sys_clk_timer_s1 OR NOT cpuNios_data_master_requests_sys_clk_timer_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_sys_clk_timer_s1 OR NOT cpuNios_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_sys_clk_timer_s1 OR NOT cpuNios_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_sysid_control_slave OR NOT cpuNios_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_sysid_control_slave OR NOT cpuNios_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_qualified_request_tse_mac_control_port OR NOT cpuNios_data_master_requests_tse_mac_control_port)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_tse_mac_control_port OR NOT ((cpuNios_data_master_read OR cpuNios_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT tse_mac_control_port_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_read OR cpuNios_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_data_master_qualified_request_tse_mac_control_port OR NOT ((cpuNios_data_master_read OR cpuNios_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT tse_mac_control_port_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_read OR cpuNios_data_master_write)))))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpuNios_data_master_address_to_slave <= cpuNios_data_master_address(26 DOWNTO 0);
  --cpuNios/data_master readdata mux, which is an e_mux
  cpuNios_data_master_readdata <= ((((((((((((((A_REP(NOT cpuNios_data_master_requests_cpuNios_jtag_debug_module, 32) OR cpuNios_jtag_debug_module_readdata_from_sa)) AND ((A_REP(NOT cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1, 32) OR registered_cpuNios_data_master_readdata))) AND ((A_REP(NOT cpuNios_data_master_requests_descriptor_memory_s1, 32) OR descriptor_memory_s1_readdata_from_sa))) AND ((A_REP(NOT cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0, 32) OR registered_cpuNios_data_master_readdata))) AND ((A_REP(NOT cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave, 32) OR registered_cpuNios_data_master_readdata))) AND ((A_REP(NOT cpuNios_data_master_requests_lcd_i2c_en_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_en_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpuNios_data_master_requests_lcd_i2c_scl_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_scl_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpuNios_data_master_requests_lcd_i2c_sdat_s1, 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_sdat_s1_readdata_from_sa)))))) AND ((A_REP(NOT cpuNios_data_master_requests_performance_counter_control_slave, 32) OR performance_counter_control_slave_readdata_from_sa))) AND ((A_REP(NOT cpuNios_data_master_requests_sgdma_rx_csr, 32) OR sgdma_rx_csr_readdata_from_sa))) AND ((A_REP(NOT cpuNios_data_master_requests_sgdma_tx_csr, 32) OR sgdma_tx_csr_readdata_from_sa))) AND ((A_REP(NOT cpuNios_data_master_requests_sys_clk_timer_s1, 32) OR (std_logic_vector'("0000000000000000") & (sys_clk_timer_s1_readdata_from_sa))))) AND ((A_REP(NOT cpuNios_data_master_requests_sysid_control_slave, 32) OR sysid_control_slave_readdata_from_sa))) AND ((A_REP(NOT cpuNios_data_master_requests_tse_mac_control_port, 32) OR registered_cpuNios_data_master_readdata));
  --actual waitrequest port, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpuNios_data_master_waitrequest <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      internal_cpuNios_data_master_waitrequest <= Vector_To_Std_Logic(NOT (A_WE_StdLogicVector((std_logic'((NOT ((cpuNios_data_master_read OR cpuNios_data_master_write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_data_master_run AND internal_cpuNios_data_master_waitrequest))))))));
    end if;

  end process;

  --unpredictable registered wait state incoming data, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      registered_cpuNios_data_master_readdata <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      registered_cpuNios_data_master_readdata <= p1_registered_cpuNios_data_master_readdata;
    end if;

  end process;

  --registered readdata mux, which is an e_mux
  p1_registered_cpuNios_data_master_readdata <= ((((A_REP(NOT cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1, 32) OR cpu_ddr_clock_bridge_s1_readdata_from_sa)) AND ((A_REP(NOT cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0, 32) OR fft_pipeline_0_avalon_slave_0_readdata_from_sa))) AND ((A_REP(NOT cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave, 32) OR jtag_uart_avalon_jtag_slave_readdata_from_sa))) AND ((A_REP(NOT cpuNios_data_master_requests_tse_mac_control_port, 32) OR tse_mac_control_port_readdata_from_sa));
  --irq assign, which is an e_assign
  cpuNios_data_master_irq <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(sys_clk_timer_s1_irq_from_sa) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(sgdma_tx_csr_irq_from_sa) & A_ToStdLogicVector(clk100MHz_lcd_sgdma_csr_irq_from_sa) & A_ToStdLogicVector(sgdma_rx_csr_irq_from_sa) & A_ToStdLogicVector(jtag_uart_avalon_jtag_slave_irq_from_sa));
  --lcd_sgdma_csr_irq_from_sa from sdram_phy_clk_out to clk100MHz
  lcd_sgdma_csr_irq_from_sa_clock_crossing_cpuNios_data_master : lcd_sgdma_csr_irq_from_sa_clock_crossing_cpuNios_data_master_module
    port map(
      data_out => clk100MHz_lcd_sgdma_csr_irq_from_sa,
      clk => clk100MHz,
      data_in => lcd_sgdma_csr_irq_from_sa,
      reset_n => clk100MHz_reset_n
    );


  --vhdl renameroo for output signals
  cpuNios_data_master_address_to_slave <= internal_cpuNios_data_master_address_to_slave;
  --vhdl renameroo for output signals
  cpuNios_data_master_waitrequest <= internal_cpuNios_data_master_waitrequest;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpuNios_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_instruction_master_address : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_instruction_master_granted_cpuNios_jtag_debug_module : IN STD_LOGIC;
                 signal cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module : IN STD_LOGIC;
                 signal cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpuNios_instruction_master_read : IN STD_LOGIC;
                 signal cpuNios_instruction_master_read_data_valid_cpuNios_jtag_debug_module : IN STD_LOGIC;
                 signal cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpuNios_instruction_master_requests_cpuNios_jtag_debug_module : IN STD_LOGIC;
                 signal cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal cpuNios_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal d1_cpuNios_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_cpu_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpuNios_instruction_master_waitrequest : OUT STD_LOGIC
              );
end entity cpuNios_instruction_master_arbitrator;


architecture europa of cpuNios_instruction_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpuNios_instruction_master_address_last_time :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal cpuNios_instruction_master_read_last_time :  STD_LOGIC;
                signal cpuNios_instruction_master_run :  STD_LOGIC;
                signal internal_cpuNios_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal internal_cpuNios_instruction_master_waitrequest :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module OR NOT cpuNios_instruction_master_requests_cpuNios_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_instruction_master_granted_cpuNios_jtag_debug_module OR NOT cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module OR NOT cpuNios_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cpuNios_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_instruction_master_read)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 OR cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1) OR NOT cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 OR NOT cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 OR NOT cpuNios_instruction_master_read) OR ((cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 AND cpuNios_instruction_master_read)))))))));
  --cascaded wait assignment, which is an e_assign
  cpuNios_instruction_master_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_cpuNios_instruction_master_address_to_slave <= cpuNios_instruction_master_address(26 DOWNTO 0);
  --cpuNios/instruction_master readdata mux, which is an e_mux
  cpuNios_instruction_master_readdata <= ((A_REP(NOT cpuNios_instruction_master_requests_cpuNios_jtag_debug_module, 32) OR cpuNios_jtag_debug_module_readdata_from_sa)) AND ((A_REP(NOT cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1, 32) OR cpu_ddr_clock_bridge_s1_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_cpuNios_instruction_master_waitrequest <= NOT cpuNios_instruction_master_run;
  --vhdl renameroo for output signals
  cpuNios_instruction_master_address_to_slave <= internal_cpuNios_instruction_master_address_to_slave;
  --vhdl renameroo for output signals
  cpuNios_instruction_master_waitrequest <= internal_cpuNios_instruction_master_waitrequest;
--synthesis translate_off
    --cpuNios_instruction_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpuNios_instruction_master_address_last_time <= std_logic_vector'("000000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpuNios_instruction_master_address_last_time <= cpuNios_instruction_master_address;
      end if;

    end process;

    --cpuNios/instruction_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpuNios_instruction_master_waitrequest AND (cpuNios_instruction_master_read);
      end if;

    end process;

    --cpuNios_instruction_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line2 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpuNios_instruction_master_address /= cpuNios_instruction_master_address_last_time))))) = '1' then 
          write(write_line2, now);
          write(write_line2, string'(": "));
          write(write_line2, string'("cpuNios_instruction_master_address did not heed wait!!!"));
          write(output, write_line2.all);
          deallocate (write_line2);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpuNios_instruction_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpuNios_instruction_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpuNios_instruction_master_read_last_time <= cpuNios_instruction_master_read;
      end if;

    end process;

    --cpuNios_instruction_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line3 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpuNios_instruction_master_read) /= std_logic'(cpuNios_instruction_master_read_last_time)))))) = '1' then 
          write(write_line3, now);
          write(write_line3, string'(": "));
          write(write_line3, string'("cpuNios_instruction_master_read did not heed wait!!!"));
          write(output, write_line3.all);
          deallocate (write_line3);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpuNios_data_master_to_cpu_ddr_clock_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpuNios_data_master_to_cpu_ddr_clock_bridge_s1_module;


architecture europa of rdv_fifo_for_cpuNios_data_master_to_cpu_ddr_clock_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_33 :  STD_LOGIC;
                signal full_34 :  STD_LOGIC;
                signal full_35 :  STD_LOGIC;
                signal full_36 :  STD_LOGIC;
                signal full_37 :  STD_LOGIC;
                signal full_38 :  STD_LOGIC;
                signal full_39 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_40 :  STD_LOGIC;
                signal full_41 :  STD_LOGIC;
                signal full_42 :  STD_LOGIC;
                signal full_43 :  STD_LOGIC;
                signal full_44 :  STD_LOGIC;
                signal full_45 :  STD_LOGIC;
                signal full_46 :  STD_LOGIC;
                signal full_47 :  STD_LOGIC;
                signal full_48 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p32_full_32 :  STD_LOGIC;
                signal p32_stage_32 :  STD_LOGIC;
                signal p33_full_33 :  STD_LOGIC;
                signal p33_stage_33 :  STD_LOGIC;
                signal p34_full_34 :  STD_LOGIC;
                signal p34_stage_34 :  STD_LOGIC;
                signal p35_full_35 :  STD_LOGIC;
                signal p35_stage_35 :  STD_LOGIC;
                signal p36_full_36 :  STD_LOGIC;
                signal p36_stage_36 :  STD_LOGIC;
                signal p37_full_37 :  STD_LOGIC;
                signal p37_stage_37 :  STD_LOGIC;
                signal p38_full_38 :  STD_LOGIC;
                signal p38_stage_38 :  STD_LOGIC;
                signal p39_full_39 :  STD_LOGIC;
                signal p39_stage_39 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p40_full_40 :  STD_LOGIC;
                signal p40_stage_40 :  STD_LOGIC;
                signal p41_full_41 :  STD_LOGIC;
                signal p41_stage_41 :  STD_LOGIC;
                signal p42_full_42 :  STD_LOGIC;
                signal p42_stage_42 :  STD_LOGIC;
                signal p43_full_43 :  STD_LOGIC;
                signal p43_stage_43 :  STD_LOGIC;
                signal p44_full_44 :  STD_LOGIC;
                signal p44_stage_44 :  STD_LOGIC;
                signal p45_full_45 :  STD_LOGIC;
                signal p45_stage_45 :  STD_LOGIC;
                signal p46_full_46 :  STD_LOGIC;
                signal p46_stage_46 :  STD_LOGIC;
                signal p47_full_47 :  STD_LOGIC;
                signal p47_stage_47 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_32 :  STD_LOGIC;
                signal stage_33 :  STD_LOGIC;
                signal stage_34 :  STD_LOGIC;
                signal stage_35 :  STD_LOGIC;
                signal stage_36 :  STD_LOGIC;
                signal stage_37 :  STD_LOGIC;
                signal stage_38 :  STD_LOGIC;
                signal stage_39 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_40 :  STD_LOGIC;
                signal stage_41 :  STD_LOGIC;
                signal stage_42 :  STD_LOGIC;
                signal stage_43 :  STD_LOGIC;
                signal stage_44 :  STD_LOGIC;
                signal stage_45 :  STD_LOGIC;
                signal stage_46 :  STD_LOGIC;
                signal stage_47 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_47;
  empty <= NOT(full_0);
  full_48 <= std_logic'('0');
  --data_47, which is an e_mux
  p47_stage_47 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_48 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_47, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_47 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_47))))) = '1' then 
        if std_logic'(((sync_reset AND full_47) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_48))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_47 <= std_logic'('0');
        else
          stage_47 <= p47_stage_47;
        end if;
      end if;
    end if;

  end process;

  --control_47, which is an e_mux
  p47_full_47 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_46))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_47, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_47 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_47 <= std_logic'('0');
        else
          full_47 <= p47_full_47;
        end if;
      end if;
    end if;

  end process;

  --data_46, which is an e_mux
  p46_stage_46 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_47 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_47);
  --data_reg_46, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_46 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_46))))) = '1' then 
        if std_logic'(((sync_reset AND full_46) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_47))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_46 <= std_logic'('0');
        else
          stage_46 <= p46_stage_46;
        end if;
      end if;
    end if;

  end process;

  --control_46, which is an e_mux
  p46_full_46 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_45, full_47);
  --control_reg_46, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_46 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_46 <= std_logic'('0');
        else
          full_46 <= p46_full_46;
        end if;
      end if;
    end if;

  end process;

  --data_45, which is an e_mux
  p45_stage_45 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_46 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_46);
  --data_reg_45, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_45 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_45))))) = '1' then 
        if std_logic'(((sync_reset AND full_45) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_46))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_45 <= std_logic'('0');
        else
          stage_45 <= p45_stage_45;
        end if;
      end if;
    end if;

  end process;

  --control_45, which is an e_mux
  p45_full_45 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_44, full_46);
  --control_reg_45, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_45 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_45 <= std_logic'('0');
        else
          full_45 <= p45_full_45;
        end if;
      end if;
    end if;

  end process;

  --data_44, which is an e_mux
  p44_stage_44 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_45 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_45);
  --data_reg_44, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_44 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_44))))) = '1' then 
        if std_logic'(((sync_reset AND full_44) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_45))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_44 <= std_logic'('0');
        else
          stage_44 <= p44_stage_44;
        end if;
      end if;
    end if;

  end process;

  --control_44, which is an e_mux
  p44_full_44 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_43, full_45);
  --control_reg_44, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_44 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_44 <= std_logic'('0');
        else
          full_44 <= p44_full_44;
        end if;
      end if;
    end if;

  end process;

  --data_43, which is an e_mux
  p43_stage_43 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_44 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_44);
  --data_reg_43, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_43 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_43))))) = '1' then 
        if std_logic'(((sync_reset AND full_43) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_44))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_43 <= std_logic'('0');
        else
          stage_43 <= p43_stage_43;
        end if;
      end if;
    end if;

  end process;

  --control_43, which is an e_mux
  p43_full_43 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_42, full_44);
  --control_reg_43, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_43 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_43 <= std_logic'('0');
        else
          full_43 <= p43_full_43;
        end if;
      end if;
    end if;

  end process;

  --data_42, which is an e_mux
  p42_stage_42 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_43 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_43);
  --data_reg_42, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_42 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_42))))) = '1' then 
        if std_logic'(((sync_reset AND full_42) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_43))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_42 <= std_logic'('0');
        else
          stage_42 <= p42_stage_42;
        end if;
      end if;
    end if;

  end process;

  --control_42, which is an e_mux
  p42_full_42 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_41, full_43);
  --control_reg_42, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_42 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_42 <= std_logic'('0');
        else
          full_42 <= p42_full_42;
        end if;
      end if;
    end if;

  end process;

  --data_41, which is an e_mux
  p41_stage_41 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_42 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_42);
  --data_reg_41, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_41 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_41))))) = '1' then 
        if std_logic'(((sync_reset AND full_41) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_42))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_41 <= std_logic'('0');
        else
          stage_41 <= p41_stage_41;
        end if;
      end if;
    end if;

  end process;

  --control_41, which is an e_mux
  p41_full_41 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_40, full_42);
  --control_reg_41, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_41 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_41 <= std_logic'('0');
        else
          full_41 <= p41_full_41;
        end if;
      end if;
    end if;

  end process;

  --data_40, which is an e_mux
  p40_stage_40 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_41 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_41);
  --data_reg_40, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_40 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_40))))) = '1' then 
        if std_logic'(((sync_reset AND full_40) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_41))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_40 <= std_logic'('0');
        else
          stage_40 <= p40_stage_40;
        end if;
      end if;
    end if;

  end process;

  --control_40, which is an e_mux
  p40_full_40 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_39, full_41);
  --control_reg_40, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_40 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_40 <= std_logic'('0');
        else
          full_40 <= p40_full_40;
        end if;
      end if;
    end if;

  end process;

  --data_39, which is an e_mux
  p39_stage_39 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_40 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_40);
  --data_reg_39, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_39 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_39))))) = '1' then 
        if std_logic'(((sync_reset AND full_39) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_40))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_39 <= std_logic'('0');
        else
          stage_39 <= p39_stage_39;
        end if;
      end if;
    end if;

  end process;

  --control_39, which is an e_mux
  p39_full_39 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_38, full_40);
  --control_reg_39, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_39 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_39 <= std_logic'('0');
        else
          full_39 <= p39_full_39;
        end if;
      end if;
    end if;

  end process;

  --data_38, which is an e_mux
  p38_stage_38 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_39 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_39);
  --data_reg_38, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_38 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_38))))) = '1' then 
        if std_logic'(((sync_reset AND full_38) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_39))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_38 <= std_logic'('0');
        else
          stage_38 <= p38_stage_38;
        end if;
      end if;
    end if;

  end process;

  --control_38, which is an e_mux
  p38_full_38 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_37, full_39);
  --control_reg_38, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_38 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_38 <= std_logic'('0');
        else
          full_38 <= p38_full_38;
        end if;
      end if;
    end if;

  end process;

  --data_37, which is an e_mux
  p37_stage_37 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_38 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_38);
  --data_reg_37, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_37 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_37))))) = '1' then 
        if std_logic'(((sync_reset AND full_37) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_38))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_37 <= std_logic'('0');
        else
          stage_37 <= p37_stage_37;
        end if;
      end if;
    end if;

  end process;

  --control_37, which is an e_mux
  p37_full_37 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_36, full_38);
  --control_reg_37, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_37 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_37 <= std_logic'('0');
        else
          full_37 <= p37_full_37;
        end if;
      end if;
    end if;

  end process;

  --data_36, which is an e_mux
  p36_stage_36 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_37 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_37);
  --data_reg_36, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_36 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_36))))) = '1' then 
        if std_logic'(((sync_reset AND full_36) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_37))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_36 <= std_logic'('0');
        else
          stage_36 <= p36_stage_36;
        end if;
      end if;
    end if;

  end process;

  --control_36, which is an e_mux
  p36_full_36 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_35, full_37);
  --control_reg_36, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_36 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_36 <= std_logic'('0');
        else
          full_36 <= p36_full_36;
        end if;
      end if;
    end if;

  end process;

  --data_35, which is an e_mux
  p35_stage_35 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_36 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_36);
  --data_reg_35, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_35 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_35))))) = '1' then 
        if std_logic'(((sync_reset AND full_35) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_36))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_35 <= std_logic'('0');
        else
          stage_35 <= p35_stage_35;
        end if;
      end if;
    end if;

  end process;

  --control_35, which is an e_mux
  p35_full_35 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_34, full_36);
  --control_reg_35, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_35 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_35 <= std_logic'('0');
        else
          full_35 <= p35_full_35;
        end if;
      end if;
    end if;

  end process;

  --data_34, which is an e_mux
  p34_stage_34 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_35 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_35);
  --data_reg_34, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_34 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_34))))) = '1' then 
        if std_logic'(((sync_reset AND full_34) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_35))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_34 <= std_logic'('0');
        else
          stage_34 <= p34_stage_34;
        end if;
      end if;
    end if;

  end process;

  --control_34, which is an e_mux
  p34_full_34 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_33, full_35);
  --control_reg_34, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_34 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_34 <= std_logic'('0');
        else
          full_34 <= p34_full_34;
        end if;
      end if;
    end if;

  end process;

  --data_33, which is an e_mux
  p33_stage_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_34 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_34);
  --data_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_33))))) = '1' then 
        if std_logic'(((sync_reset AND full_33) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_34))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_33 <= std_logic'('0');
        else
          stage_33 <= p33_stage_33;
        end if;
      end if;
    end if;

  end process;

  --control_33, which is an e_mux
  p33_full_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_32, full_34);
  --control_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_33 <= std_logic'('0');
        else
          full_33 <= p33_full_33;
        end if;
      end if;
    end if;

  end process;

  --data_32, which is an e_mux
  p32_stage_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_33 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_33);
  --data_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_32))))) = '1' then 
        if std_logic'(((sync_reset AND full_32) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_33))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_32 <= std_logic'('0');
        else
          stage_32 <= p32_stage_32;
        end if;
      end if;
    end if;

  end process;

  --control_32, which is an e_mux
  p32_full_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_31, full_33);
  --control_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_32 <= std_logic'('0');
        else
          full_32 <= p32_full_32;
        end if;
      end if;
    end if;

  end process;

  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_32);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_30, full_32);
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpuNios_instruction_master_to_cpu_ddr_clock_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpuNios_instruction_master_to_cpu_ddr_clock_bridge_s1_module;


architecture europa of rdv_fifo_for_cpuNios_instruction_master_to_cpu_ddr_clock_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_33 :  STD_LOGIC;
                signal full_34 :  STD_LOGIC;
                signal full_35 :  STD_LOGIC;
                signal full_36 :  STD_LOGIC;
                signal full_37 :  STD_LOGIC;
                signal full_38 :  STD_LOGIC;
                signal full_39 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_40 :  STD_LOGIC;
                signal full_41 :  STD_LOGIC;
                signal full_42 :  STD_LOGIC;
                signal full_43 :  STD_LOGIC;
                signal full_44 :  STD_LOGIC;
                signal full_45 :  STD_LOGIC;
                signal full_46 :  STD_LOGIC;
                signal full_47 :  STD_LOGIC;
                signal full_48 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p32_full_32 :  STD_LOGIC;
                signal p32_stage_32 :  STD_LOGIC;
                signal p33_full_33 :  STD_LOGIC;
                signal p33_stage_33 :  STD_LOGIC;
                signal p34_full_34 :  STD_LOGIC;
                signal p34_stage_34 :  STD_LOGIC;
                signal p35_full_35 :  STD_LOGIC;
                signal p35_stage_35 :  STD_LOGIC;
                signal p36_full_36 :  STD_LOGIC;
                signal p36_stage_36 :  STD_LOGIC;
                signal p37_full_37 :  STD_LOGIC;
                signal p37_stage_37 :  STD_LOGIC;
                signal p38_full_38 :  STD_LOGIC;
                signal p38_stage_38 :  STD_LOGIC;
                signal p39_full_39 :  STD_LOGIC;
                signal p39_stage_39 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p40_full_40 :  STD_LOGIC;
                signal p40_stage_40 :  STD_LOGIC;
                signal p41_full_41 :  STD_LOGIC;
                signal p41_stage_41 :  STD_LOGIC;
                signal p42_full_42 :  STD_LOGIC;
                signal p42_stage_42 :  STD_LOGIC;
                signal p43_full_43 :  STD_LOGIC;
                signal p43_stage_43 :  STD_LOGIC;
                signal p44_full_44 :  STD_LOGIC;
                signal p44_stage_44 :  STD_LOGIC;
                signal p45_full_45 :  STD_LOGIC;
                signal p45_stage_45 :  STD_LOGIC;
                signal p46_full_46 :  STD_LOGIC;
                signal p46_stage_46 :  STD_LOGIC;
                signal p47_full_47 :  STD_LOGIC;
                signal p47_stage_47 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_32 :  STD_LOGIC;
                signal stage_33 :  STD_LOGIC;
                signal stage_34 :  STD_LOGIC;
                signal stage_35 :  STD_LOGIC;
                signal stage_36 :  STD_LOGIC;
                signal stage_37 :  STD_LOGIC;
                signal stage_38 :  STD_LOGIC;
                signal stage_39 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_40 :  STD_LOGIC;
                signal stage_41 :  STD_LOGIC;
                signal stage_42 :  STD_LOGIC;
                signal stage_43 :  STD_LOGIC;
                signal stage_44 :  STD_LOGIC;
                signal stage_45 :  STD_LOGIC;
                signal stage_46 :  STD_LOGIC;
                signal stage_47 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_47;
  empty <= NOT(full_0);
  full_48 <= std_logic'('0');
  --data_47, which is an e_mux
  p47_stage_47 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_48 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_47, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_47 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_47))))) = '1' then 
        if std_logic'(((sync_reset AND full_47) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_48))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_47 <= std_logic'('0');
        else
          stage_47 <= p47_stage_47;
        end if;
      end if;
    end if;

  end process;

  --control_47, which is an e_mux
  p47_full_47 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_46))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_47, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_47 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_47 <= std_logic'('0');
        else
          full_47 <= p47_full_47;
        end if;
      end if;
    end if;

  end process;

  --data_46, which is an e_mux
  p46_stage_46 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_47 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_47);
  --data_reg_46, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_46 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_46))))) = '1' then 
        if std_logic'(((sync_reset AND full_46) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_47))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_46 <= std_logic'('0');
        else
          stage_46 <= p46_stage_46;
        end if;
      end if;
    end if;

  end process;

  --control_46, which is an e_mux
  p46_full_46 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_45, full_47);
  --control_reg_46, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_46 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_46 <= std_logic'('0');
        else
          full_46 <= p46_full_46;
        end if;
      end if;
    end if;

  end process;

  --data_45, which is an e_mux
  p45_stage_45 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_46 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_46);
  --data_reg_45, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_45 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_45))))) = '1' then 
        if std_logic'(((sync_reset AND full_45) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_46))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_45 <= std_logic'('0');
        else
          stage_45 <= p45_stage_45;
        end if;
      end if;
    end if;

  end process;

  --control_45, which is an e_mux
  p45_full_45 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_44, full_46);
  --control_reg_45, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_45 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_45 <= std_logic'('0');
        else
          full_45 <= p45_full_45;
        end if;
      end if;
    end if;

  end process;

  --data_44, which is an e_mux
  p44_stage_44 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_45 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_45);
  --data_reg_44, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_44 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_44))))) = '1' then 
        if std_logic'(((sync_reset AND full_44) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_45))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_44 <= std_logic'('0');
        else
          stage_44 <= p44_stage_44;
        end if;
      end if;
    end if;

  end process;

  --control_44, which is an e_mux
  p44_full_44 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_43, full_45);
  --control_reg_44, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_44 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_44 <= std_logic'('0');
        else
          full_44 <= p44_full_44;
        end if;
      end if;
    end if;

  end process;

  --data_43, which is an e_mux
  p43_stage_43 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_44 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_44);
  --data_reg_43, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_43 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_43))))) = '1' then 
        if std_logic'(((sync_reset AND full_43) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_44))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_43 <= std_logic'('0');
        else
          stage_43 <= p43_stage_43;
        end if;
      end if;
    end if;

  end process;

  --control_43, which is an e_mux
  p43_full_43 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_42, full_44);
  --control_reg_43, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_43 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_43 <= std_logic'('0');
        else
          full_43 <= p43_full_43;
        end if;
      end if;
    end if;

  end process;

  --data_42, which is an e_mux
  p42_stage_42 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_43 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_43);
  --data_reg_42, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_42 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_42))))) = '1' then 
        if std_logic'(((sync_reset AND full_42) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_43))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_42 <= std_logic'('0');
        else
          stage_42 <= p42_stage_42;
        end if;
      end if;
    end if;

  end process;

  --control_42, which is an e_mux
  p42_full_42 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_41, full_43);
  --control_reg_42, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_42 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_42 <= std_logic'('0');
        else
          full_42 <= p42_full_42;
        end if;
      end if;
    end if;

  end process;

  --data_41, which is an e_mux
  p41_stage_41 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_42 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_42);
  --data_reg_41, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_41 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_41))))) = '1' then 
        if std_logic'(((sync_reset AND full_41) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_42))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_41 <= std_logic'('0');
        else
          stage_41 <= p41_stage_41;
        end if;
      end if;
    end if;

  end process;

  --control_41, which is an e_mux
  p41_full_41 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_40, full_42);
  --control_reg_41, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_41 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_41 <= std_logic'('0');
        else
          full_41 <= p41_full_41;
        end if;
      end if;
    end if;

  end process;

  --data_40, which is an e_mux
  p40_stage_40 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_41 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_41);
  --data_reg_40, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_40 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_40))))) = '1' then 
        if std_logic'(((sync_reset AND full_40) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_41))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_40 <= std_logic'('0');
        else
          stage_40 <= p40_stage_40;
        end if;
      end if;
    end if;

  end process;

  --control_40, which is an e_mux
  p40_full_40 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_39, full_41);
  --control_reg_40, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_40 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_40 <= std_logic'('0');
        else
          full_40 <= p40_full_40;
        end if;
      end if;
    end if;

  end process;

  --data_39, which is an e_mux
  p39_stage_39 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_40 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_40);
  --data_reg_39, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_39 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_39))))) = '1' then 
        if std_logic'(((sync_reset AND full_39) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_40))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_39 <= std_logic'('0');
        else
          stage_39 <= p39_stage_39;
        end if;
      end if;
    end if;

  end process;

  --control_39, which is an e_mux
  p39_full_39 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_38, full_40);
  --control_reg_39, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_39 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_39 <= std_logic'('0');
        else
          full_39 <= p39_full_39;
        end if;
      end if;
    end if;

  end process;

  --data_38, which is an e_mux
  p38_stage_38 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_39 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_39);
  --data_reg_38, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_38 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_38))))) = '1' then 
        if std_logic'(((sync_reset AND full_38) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_39))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_38 <= std_logic'('0');
        else
          stage_38 <= p38_stage_38;
        end if;
      end if;
    end if;

  end process;

  --control_38, which is an e_mux
  p38_full_38 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_37, full_39);
  --control_reg_38, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_38 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_38 <= std_logic'('0');
        else
          full_38 <= p38_full_38;
        end if;
      end if;
    end if;

  end process;

  --data_37, which is an e_mux
  p37_stage_37 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_38 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_38);
  --data_reg_37, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_37 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_37))))) = '1' then 
        if std_logic'(((sync_reset AND full_37) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_38))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_37 <= std_logic'('0');
        else
          stage_37 <= p37_stage_37;
        end if;
      end if;
    end if;

  end process;

  --control_37, which is an e_mux
  p37_full_37 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_36, full_38);
  --control_reg_37, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_37 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_37 <= std_logic'('0');
        else
          full_37 <= p37_full_37;
        end if;
      end if;
    end if;

  end process;

  --data_36, which is an e_mux
  p36_stage_36 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_37 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_37);
  --data_reg_36, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_36 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_36))))) = '1' then 
        if std_logic'(((sync_reset AND full_36) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_37))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_36 <= std_logic'('0');
        else
          stage_36 <= p36_stage_36;
        end if;
      end if;
    end if;

  end process;

  --control_36, which is an e_mux
  p36_full_36 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_35, full_37);
  --control_reg_36, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_36 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_36 <= std_logic'('0');
        else
          full_36 <= p36_full_36;
        end if;
      end if;
    end if;

  end process;

  --data_35, which is an e_mux
  p35_stage_35 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_36 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_36);
  --data_reg_35, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_35 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_35))))) = '1' then 
        if std_logic'(((sync_reset AND full_35) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_36))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_35 <= std_logic'('0');
        else
          stage_35 <= p35_stage_35;
        end if;
      end if;
    end if;

  end process;

  --control_35, which is an e_mux
  p35_full_35 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_34, full_36);
  --control_reg_35, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_35 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_35 <= std_logic'('0');
        else
          full_35 <= p35_full_35;
        end if;
      end if;
    end if;

  end process;

  --data_34, which is an e_mux
  p34_stage_34 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_35 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_35);
  --data_reg_34, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_34 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_34))))) = '1' then 
        if std_logic'(((sync_reset AND full_34) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_35))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_34 <= std_logic'('0');
        else
          stage_34 <= p34_stage_34;
        end if;
      end if;
    end if;

  end process;

  --control_34, which is an e_mux
  p34_full_34 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_33, full_35);
  --control_reg_34, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_34 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_34 <= std_logic'('0');
        else
          full_34 <= p34_full_34;
        end if;
      end if;
    end if;

  end process;

  --data_33, which is an e_mux
  p33_stage_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_34 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_34);
  --data_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_33))))) = '1' then 
        if std_logic'(((sync_reset AND full_33) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_34))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_33 <= std_logic'('0');
        else
          stage_33 <= p33_stage_33;
        end if;
      end if;
    end if;

  end process;

  --control_33, which is an e_mux
  p33_full_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_32, full_34);
  --control_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_33 <= std_logic'('0');
        else
          full_33 <= p33_full_33;
        end if;
      end if;
    end if;

  end process;

  --data_32, which is an e_mux
  p32_stage_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_33 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_33);
  --data_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_32))))) = '1' then 
        if std_logic'(((sync_reset AND full_32) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_33))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_32 <= std_logic'('0');
        else
          stage_32 <= p32_stage_32;
        end if;
      end if;
    end if;

  end process;

  --control_32, which is an e_mux
  p32_full_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_31, full_33);
  --control_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_32 <= std_logic'('0');
        else
          full_32 <= p32_full_32;
        end if;
      end if;
    end if;

  end process;

  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_32);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_30, full_32);
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_ddr_clock_bridge_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpuNios_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_instruction_master_read : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_endofpacket : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_readdatavalid : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_read : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_s1_reset_n : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_write : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_ddr_clock_bridge_s1_end_xfer : OUT STD_LOGIC
              );
end entity cpu_ddr_clock_bridge_s1_arbitrator;


architecture europa of cpu_ddr_clock_bridge_s1_arbitrator is
component rdv_fifo_for_cpuNios_data_master_to_cpu_ddr_clock_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpuNios_data_master_to_cpu_ddr_clock_bridge_s1_module;

component rdv_fifo_for_cpuNios_instruction_master_to_cpu_ddr_clock_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpuNios_instruction_master_to_cpu_ddr_clock_bridge_s1_module;

                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_data_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_instruction_master_continuerequest :  STD_LOGIC;
                signal cpuNios_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_instruction_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_allgrants :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_any_continuerequest :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_arb_counter_enable :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_begins_xfer :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_end_xfer :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_firsttransfer :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_in_a_read_cycle :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_in_a_write_cycle :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_non_bursting_master_requests :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_reg_firsttransfer :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_slavearbiterlockenable :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_unreg_firsttransfer :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_waits_for_read :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register :  STD_LOGIC;
                signal internal_cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_cpuNios_data_master_granted_slave_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal last_cycle_cpuNios_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal module_input :  STD_LOGIC;
                signal module_input1 :  STD_LOGIC;
                signal module_input2 :  STD_LOGIC;
                signal module_input3 :  STD_LOGIC;
                signal module_input4 :  STD_LOGIC;
                signal module_input5 :  STD_LOGIC;
                signal shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpuNios_instruction_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_cpu_ddr_clock_bridge_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cpu_ddr_clock_bridge_s1_end_xfer;
    end if;

  end process;

  cpu_ddr_clock_bridge_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 OR internal_cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1));
  --assign cpu_ddr_clock_bridge_s1_readdata_from_sa = cpu_ddr_clock_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_ddr_clock_bridge_s1_readdata_from_sa <= cpu_ddr_clock_bridge_s1_readdata;
  internal_cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 <= to_std_logic(((Std_Logic_Vector'(A_ToStdLogicVector(cpuNios_data_master_address_to_slave(26)) & std_logic_vector'("00000000000000000000000000")) = std_logic_vector'("000000000000000000000000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --assign cpu_ddr_clock_bridge_s1_waitrequest_from_sa = cpu_ddr_clock_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_cpu_ddr_clock_bridge_s1_waitrequest_from_sa <= cpu_ddr_clock_bridge_s1_waitrequest;
  --assign cpu_ddr_clock_bridge_s1_readdatavalid_from_sa = cpu_ddr_clock_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_ddr_clock_bridge_s1_readdatavalid_from_sa <= cpu_ddr_clock_bridge_s1_readdatavalid;
  --cpu_ddr_clock_bridge_s1_arb_share_counter set values, which is an e_mux
  cpu_ddr_clock_bridge_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), std_logic_vector'("00000000000000000000000000000001"))))), 4);
  --cpu_ddr_clock_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_non_bursting_master_requests <= ((internal_cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 OR internal_cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1) OR internal_cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1) OR internal_cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  --cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --cpu_ddr_clock_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  cpu_ddr_clock_bridge_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(cpu_ddr_clock_bridge_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (cpu_ddr_clock_bridge_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(cpu_ddr_clock_bridge_s1_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (cpu_ddr_clock_bridge_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --cpu_ddr_clock_bridge_s1_allgrants all slave grants, which is an e_mux
  cpu_ddr_clock_bridge_s1_allgrants <= (((or_reduce(cpu_ddr_clock_bridge_s1_grant_vector)) OR (or_reduce(cpu_ddr_clock_bridge_s1_grant_vector))) OR (or_reduce(cpu_ddr_clock_bridge_s1_grant_vector))) OR (or_reduce(cpu_ddr_clock_bridge_s1_grant_vector));
  --cpu_ddr_clock_bridge_s1_end_xfer assignment, which is an e_assign
  cpu_ddr_clock_bridge_s1_end_xfer <= NOT ((cpu_ddr_clock_bridge_s1_waits_for_read OR cpu_ddr_clock_bridge_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 <= cpu_ddr_clock_bridge_s1_end_xfer AND (((NOT cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cpu_ddr_clock_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  cpu_ddr_clock_bridge_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 AND cpu_ddr_clock_bridge_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 AND NOT cpu_ddr_clock_bridge_s1_non_bursting_master_requests));
  --cpu_ddr_clock_bridge_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_s1_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_ddr_clock_bridge_s1_arb_counter_enable) = '1' then 
        cpu_ddr_clock_bridge_s1_arb_share_counter <= cpu_ddr_clock_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_ddr_clock_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(cpu_ddr_clock_bridge_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1)) OR ((end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 AND NOT cpu_ddr_clock_bridge_s1_non_bursting_master_requests)))) = '1' then 
        cpu_ddr_clock_bridge_s1_slavearbiterlockenable <= or_reduce(cpu_ddr_clock_bridge_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpuNios/data_master cpu_ddr_clock_bridge/s1 arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= cpu_ddr_clock_bridge_s1_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 <= or_reduce(cpu_ddr_clock_bridge_s1_arb_share_counter_next_value);
  --cpuNios/data_master cpu_ddr_clock_bridge/s1 arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --cpuNios/instruction_master cpu_ddr_clock_bridge/s1 arbiterlock, which is an e_assign
  cpuNios_instruction_master_arbiterlock <= cpu_ddr_clock_bridge_s1_slavearbiterlockenable AND cpuNios_instruction_master_continuerequest;
  --cpuNios/instruction_master cpu_ddr_clock_bridge/s1 arbiterlock2, which is an e_assign
  cpuNios_instruction_master_arbiterlock2 <= cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 AND cpuNios_instruction_master_continuerequest;
  --cpuNios/instruction_master granted cpu_ddr_clock_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpuNios_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpuNios_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpuNios_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal OR NOT internal_cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpuNios_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1))))));
    end if;

  end process;

  --cpuNios_instruction_master_continuerequest continued request, which is an e_mux
  cpuNios_instruction_master_continuerequest <= last_cycle_cpuNios_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 AND internal_cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  --cpu_ddr_clock_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  cpu_ddr_clock_bridge_s1_any_continuerequest <= cpuNios_instruction_master_continuerequest OR cpuNios_data_master_continuerequest;
  internal_cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 <= internal_cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 AND NOT (((((cpuNios_data_master_read AND ((NOT cpuNios_data_master_waitrequest OR (internal_cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register))))) OR (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write))) OR cpuNios_instruction_master_arbiterlock));
  --unique name for cpu_ddr_clock_bridge_s1_move_on_to_next_transaction, which is an e_assign
  cpu_ddr_clock_bridge_s1_move_on_to_next_transaction <= cpu_ddr_clock_bridge_s1_readdatavalid_from_sa;
  --rdv_fifo_for_cpuNios_data_master_to_cpu_ddr_clock_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpuNios_data_master_to_cpu_ddr_clock_bridge_s1 : rdv_fifo_for_cpuNios_data_master_to_cpu_ddr_clock_bridge_s1_module
    port map(
      data_out => cpuNios_data_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1,
      empty => open,
      fifo_contains_ones_n => cpuNios_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1,
      full => open,
      clear_fifo => module_input,
      clk => clk,
      data_in => internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1,
      read => cpu_ddr_clock_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input1,
      write => module_input2
    );

  module_input <= std_logic'('0');
  module_input1 <= std_logic'('0');
  module_input2 <= in_a_read_cycle AND NOT cpu_ddr_clock_bridge_s1_waits_for_read;

  internal_cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register <= NOT cpuNios_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  --local readdatavalid cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1, which is an e_mux
  cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 <= ((cpu_ddr_clock_bridge_s1_readdatavalid_from_sa AND cpuNios_data_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1)) AND NOT cpuNios_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  --cpu_ddr_clock_bridge_s1_writedata mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_writedata <= cpuNios_data_master_writedata;
  --assign cpu_ddr_clock_bridge_s1_endofpacket_from_sa = cpu_ddr_clock_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_ddr_clock_bridge_s1_endofpacket_from_sa <= cpu_ddr_clock_bridge_s1_endofpacket;
  internal_cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 <= ((to_std_logic(((Std_Logic_Vector'(A_ToStdLogicVector(cpuNios_instruction_master_address_to_slave(26)) & std_logic_vector'("00000000000000000000000000")) = std_logic_vector'("000000000000000000000000000")))) AND (cpuNios_instruction_master_read))) AND cpuNios_instruction_master_read;
  --cpuNios/data_master granted cpu_ddr_clock_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpuNios_data_master_granted_slave_cpu_ddr_clock_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpuNios_data_master_granted_slave_cpu_ddr_clock_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpuNios_data_master_saved_grant_cpu_ddr_clock_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal OR NOT internal_cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpuNios_data_master_granted_slave_cpu_ddr_clock_bridge_s1))))));
    end if;

  end process;

  --cpuNios_data_master_continuerequest continued request, which is an e_mux
  cpuNios_data_master_continuerequest <= last_cycle_cpuNios_data_master_granted_slave_cpu_ddr_clock_bridge_s1 AND internal_cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1;
  internal_cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 <= internal_cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 AND NOT ((((cpuNios_instruction_master_read AND (internal_cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register))) OR cpuNios_data_master_arbiterlock));
  --rdv_fifo_for_cpuNios_instruction_master_to_cpu_ddr_clock_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpuNios_instruction_master_to_cpu_ddr_clock_bridge_s1 : rdv_fifo_for_cpuNios_instruction_master_to_cpu_ddr_clock_bridge_s1_module
    port map(
      data_out => cpuNios_instruction_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1,
      empty => open,
      fifo_contains_ones_n => cpuNios_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1,
      full => open,
      clear_fifo => module_input3,
      clk => clk,
      data_in => internal_cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1,
      read => cpu_ddr_clock_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input4,
      write => module_input5
    );

  module_input3 <= std_logic'('0');
  module_input4 <= std_logic'('0');
  module_input5 <= in_a_read_cycle AND NOT cpu_ddr_clock_bridge_s1_waits_for_read;

  internal_cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register <= NOT cpuNios_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  --local readdatavalid cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1, which is an e_mux
  cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 <= ((cpu_ddr_clock_bridge_s1_readdatavalid_from_sa AND cpuNios_instruction_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1)) AND NOT cpuNios_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  --allow new arb cycle for cpu_ddr_clock_bridge/s1, which is an e_assign
  cpu_ddr_clock_bridge_s1_allow_new_arb_cycle <= NOT cpuNios_data_master_arbiterlock AND NOT cpuNios_instruction_master_arbiterlock;
  --cpuNios/instruction_master assignment into master qualified-requests vector for cpu_ddr_clock_bridge/s1, which is an e_assign
  cpu_ddr_clock_bridge_s1_master_qreq_vector(0) <= internal_cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1;
  --cpuNios/instruction_master grant cpu_ddr_clock_bridge/s1, which is an e_assign
  internal_cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 <= cpu_ddr_clock_bridge_s1_grant_vector(0);
  --cpuNios/instruction_master saved-grant cpu_ddr_clock_bridge/s1, which is an e_assign
  cpuNios_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1 <= cpu_ddr_clock_bridge_s1_arb_winner(0) AND internal_cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  --cpuNios/data_master assignment into master qualified-requests vector for cpu_ddr_clock_bridge/s1, which is an e_assign
  cpu_ddr_clock_bridge_s1_master_qreq_vector(1) <= internal_cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1;
  --cpuNios/data_master grant cpu_ddr_clock_bridge/s1, which is an e_assign
  internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 <= cpu_ddr_clock_bridge_s1_grant_vector(1);
  --cpuNios/data_master saved-grant cpu_ddr_clock_bridge/s1, which is an e_assign
  cpuNios_data_master_saved_grant_cpu_ddr_clock_bridge_s1 <= cpu_ddr_clock_bridge_s1_arb_winner(1) AND internal_cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1;
  --cpu_ddr_clock_bridge/s1 chosen-master double-vector, which is an e_assign
  cpu_ddr_clock_bridge_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((cpu_ddr_clock_bridge_s1_master_qreq_vector & cpu_ddr_clock_bridge_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT cpu_ddr_clock_bridge_s1_master_qreq_vector & NOT cpu_ddr_clock_bridge_s1_master_qreq_vector))) + (std_logic_vector'("000") & (cpu_ddr_clock_bridge_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  cpu_ddr_clock_bridge_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((cpu_ddr_clock_bridge_s1_allow_new_arb_cycle AND or_reduce(cpu_ddr_clock_bridge_s1_grant_vector)))) = '1'), cpu_ddr_clock_bridge_s1_grant_vector, cpu_ddr_clock_bridge_s1_saved_chosen_master_vector);
  --saved cpu_ddr_clock_bridge_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_ddr_clock_bridge_s1_allow_new_arb_cycle) = '1' then 
        cpu_ddr_clock_bridge_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(cpu_ddr_clock_bridge_s1_grant_vector)) = '1'), cpu_ddr_clock_bridge_s1_grant_vector, cpu_ddr_clock_bridge_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  cpu_ddr_clock_bridge_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((cpu_ddr_clock_bridge_s1_chosen_master_double_vector(1) OR cpu_ddr_clock_bridge_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((cpu_ddr_clock_bridge_s1_chosen_master_double_vector(0) OR cpu_ddr_clock_bridge_s1_chosen_master_double_vector(2)))));
  --cpu_ddr_clock_bridge/s1 chosen master rotated left, which is an e_assign
  cpu_ddr_clock_bridge_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(cpu_ddr_clock_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(cpu_ddr_clock_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --cpu_ddr_clock_bridge/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(cpu_ddr_clock_bridge_s1_grant_vector)) = '1' then 
        cpu_ddr_clock_bridge_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(cpu_ddr_clock_bridge_s1_end_xfer) = '1'), cpu_ddr_clock_bridge_s1_chosen_master_rot_left, cpu_ddr_clock_bridge_s1_grant_vector);
      end if;
    end if;

  end process;

  --cpu_ddr_clock_bridge_s1_reset_n assignment, which is an e_assign
  cpu_ddr_clock_bridge_s1_reset_n <= reset_n;
  --cpu_ddr_clock_bridge_s1_firsttransfer first transaction, which is an e_assign
  cpu_ddr_clock_bridge_s1_firsttransfer <= A_WE_StdLogic((std_logic'(cpu_ddr_clock_bridge_s1_begins_xfer) = '1'), cpu_ddr_clock_bridge_s1_unreg_firsttransfer, cpu_ddr_clock_bridge_s1_reg_firsttransfer);
  --cpu_ddr_clock_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  cpu_ddr_clock_bridge_s1_unreg_firsttransfer <= NOT ((cpu_ddr_clock_bridge_s1_slavearbiterlockenable AND cpu_ddr_clock_bridge_s1_any_continuerequest));
  --cpu_ddr_clock_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_ddr_clock_bridge_s1_begins_xfer) = '1' then 
        cpu_ddr_clock_bridge_s1_reg_firsttransfer <= cpu_ddr_clock_bridge_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cpu_ddr_clock_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cpu_ddr_clock_bridge_s1_beginbursttransfer_internal <= cpu_ddr_clock_bridge_s1_begins_xfer;
  --cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal <= cpu_ddr_clock_bridge_s1_begins_xfer AND cpu_ddr_clock_bridge_s1_firsttransfer;
  --cpu_ddr_clock_bridge_s1_read assignment, which is an e_mux
  cpu_ddr_clock_bridge_s1_read <= ((internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 AND cpuNios_data_master_read)) OR ((internal_cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 AND cpuNios_instruction_master_read));
  --cpu_ddr_clock_bridge_s1_write assignment, which is an e_mux
  cpu_ddr_clock_bridge_s1_write <= internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 AND cpuNios_data_master_write;
  shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --cpu_ddr_clock_bridge_s1_address mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1)) = '1'), (A_SRL(shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpuNios_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 24);
  shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpuNios_instruction_master <= cpuNios_instruction_master_address_to_slave;
  --slaveid cpu_ddr_clock_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_nativeaddress <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1)) = '1'), (A_SRL(cpuNios_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(cpuNios_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")))), 24);
  --d1_cpu_ddr_clock_bridge_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cpu_ddr_clock_bridge_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cpu_ddr_clock_bridge_s1_end_xfer <= cpu_ddr_clock_bridge_s1_end_xfer;
    end if;

  end process;

  --cpu_ddr_clock_bridge_s1_waits_for_read in a cycle, which is an e_mux
  cpu_ddr_clock_bridge_s1_waits_for_read <= cpu_ddr_clock_bridge_s1_in_a_read_cycle AND internal_cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  --cpu_ddr_clock_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  cpu_ddr_clock_bridge_s1_in_a_read_cycle <= ((internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 AND cpuNios_data_master_read)) OR ((internal_cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 AND cpuNios_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cpu_ddr_clock_bridge_s1_in_a_read_cycle;
  --cpu_ddr_clock_bridge_s1_waits_for_write in a cycle, which is an e_mux
  cpu_ddr_clock_bridge_s1_waits_for_write <= cpu_ddr_clock_bridge_s1_in_a_write_cycle AND internal_cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  --cpu_ddr_clock_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  cpu_ddr_clock_bridge_s1_in_a_write_cycle <= internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cpu_ddr_clock_bridge_s1_in_a_write_cycle;
  wait_for_cpu_ddr_clock_bridge_s1_counter <= std_logic'('0');
  --cpu_ddr_clock_bridge_s1_byteenable byte enable port mux, which is an e_mux
  cpu_ddr_clock_bridge_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpuNios_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 <= internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 <= internal_cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register <= internal_cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 <= internal_cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 <= internal_cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 <= internal_cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register <= internal_cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  --vhdl renameroo for output signals
  cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 <= internal_cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_s1_waitrequest_from_sa <= internal_cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
--synthesis translate_off
    --cpu_ddr_clock_bridge/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line4 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line4, now);
          write(write_line4, string'(": "));
          write(write_line4, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line4.all);
          deallocate (write_line4);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line5 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_saved_grant_cpu_ddr_clock_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpuNios_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line5, now);
          write(write_line5, string'(": "));
          write(write_line5, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line5.all);
          deallocate (write_line5);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_module;


architecture europa of selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_ddr_clock_bridge_m1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_granted_sdram_s1 : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_requests_sdram_s1 : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_lcd_sgdma_csr_end_xfer : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal lcd_sgdma_csr_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal cpu_ddr_clock_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_latency_counter : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_readdatavalid : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_reset_n : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_waitrequest : OUT STD_LOGIC
              );
end entity cpu_ddr_clock_bridge_m1_arbitrator;


architecture europa of cpu_ddr_clock_bridge_m1_arbitrator is
component selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_module;

                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_address_last_time :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_is_granted_some_slave :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_read_but_no_slave_selected :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_read_last_time :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_run :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_write_last_time :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal empty_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo :  STD_LOGIC;
                signal full_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal internal_cpu_ddr_clock_bridge_m1_latency_counter :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal module_input6 :  STD_LOGIC;
                signal module_input7 :  STD_LOGIC;
                signal module_input8 :  STD_LOGIC;
                signal p1_cpu_ddr_clock_bridge_m1_latency_counter :  STD_LOGIC;
                signal pre_flush_cpu_ddr_clock_bridge_m1_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal read_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo :  STD_LOGIC;
                signal sdram_s1_readdata_from_sa_part_selected_by_negative_dbs :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_output :  STD_LOGIC;
                signal selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_output_sdram_s1 :  STD_LOGIC;
                signal write_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr OR NOT cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr OR NOT cpu_ddr_clock_bridge_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_lcd_sgdma_csr_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr OR NOT cpu_ddr_clock_bridge_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 OR NOT cpu_ddr_clock_bridge_m1_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_ddr_clock_bridge_m1_granted_sdram_s1 OR NOT cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 OR NOT ((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 OR NOT ((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_ddr_clock_bridge_m1_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_ddr_clock_bridge_m1_address_to_slave <= cpu_ddr_clock_bridge_m1_address(25 DOWNTO 0);
  --cpu_ddr_clock_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_ddr_clock_bridge_m1_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_ddr_clock_bridge_m1_read_but_no_slave_selected <= (cpu_ddr_clock_bridge_m1_read AND cpu_ddr_clock_bridge_m1_run) AND NOT cpu_ddr_clock_bridge_m1_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  cpu_ddr_clock_bridge_m1_is_granted_some_slave <= cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr OR cpu_ddr_clock_bridge_m1_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_cpu_ddr_clock_bridge_m1_readdatavalid <= cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  cpu_ddr_clock_bridge_m1_readdatavalid <= (((cpu_ddr_clock_bridge_m1_read_but_no_slave_selected OR pre_flush_cpu_ddr_clock_bridge_m1_readdatavalid) OR cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr) OR cpu_ddr_clock_bridge_m1_read_but_no_slave_selected) OR pre_flush_cpu_ddr_clock_bridge_m1_readdatavalid;
  --cpu_ddr_clock_bridge/m1 readdata mux, which is an e_mux
  cpu_ddr_clock_bridge_m1_readdata <= ((A_REP(NOT ((cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr AND cpu_ddr_clock_bridge_m1_read)) , 32) OR lcd_sgdma_csr_readdata_from_sa)) AND ((A_REP(NOT cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1, 32) OR sdram_s1_readdata_from_sa_part_selected_by_negative_dbs));
  --actual waitrequest port, which is an e_assign
  internal_cpu_ddr_clock_bridge_m1_waitrequest <= NOT cpu_ddr_clock_bridge_m1_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_ddr_clock_bridge_m1_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_cpu_ddr_clock_bridge_m1_latency_counter <= p1_cpu_ddr_clock_bridge_m1_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_cpu_ddr_clock_bridge_m1_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((cpu_ddr_clock_bridge_m1_run AND cpu_ddr_clock_bridge_m1_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_cpu_ddr_clock_bridge_m1_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_cpu_ddr_clock_bridge_m1_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --cpu_ddr_clock_bridge_m1_reset_n assignment, which is an e_assign
  cpu_ddr_clock_bridge_m1_reset_n <= reset_n;
  --Negative Dynamic Bus-sizing mux.
  --this mux selects the correct half of the 
  --wide data coming from the slave sdram/s1 
  sdram_s1_readdata_from_sa_part_selected_by_negative_dbs <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_output_sdram_s1))) = std_logic_vector'("00000000000000000000000000000000"))), sdram_s1_readdata_from_sa(31 DOWNTO 0), sdram_s1_readdata_from_sa(63 DOWNTO 32));
  --read_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo fifo read, which is an e_mux
  read_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo <= cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1;
  --write_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo fifo write, which is an e_mux
  write_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo <= (cpu_ddr_clock_bridge_m1_read AND cpu_ddr_clock_bridge_m1_run) AND cpu_ddr_clock_bridge_m1_requests_sdram_s1;
  selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_output_sdram_s1 <= selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_output;
  --selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo, which is an e_fifo_with_registered_outputs
  selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo : selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_module
    port map(
      data_out => selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo_output,
      empty => empty_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo,
      fifo_contains_ones_n => open,
      full => full_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo,
      clear_fifo => module_input6,
      clk => clk,
      data_in => module_input7,
      read => read_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo,
      reset_n => reset_n,
      sync_reset => module_input8,
      write => write_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo
    );

  module_input6 <= std_logic'('0');
  module_input7 <= internal_cpu_ddr_clock_bridge_m1_address_to_slave(2);
  module_input8 <= std_logic'('0');

  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_address_to_slave <= internal_cpu_ddr_clock_bridge_m1_address_to_slave;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_latency_counter <= internal_cpu_ddr_clock_bridge_m1_latency_counter;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_waitrequest <= internal_cpu_ddr_clock_bridge_m1_waitrequest;
--synthesis translate_off
    --cpu_ddr_clock_bridge_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_ddr_clock_bridge_m1_address_last_time <= std_logic_vector'("00000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_ddr_clock_bridge_m1_address_last_time <= cpu_ddr_clock_bridge_m1_address;
      end if;

    end process;

    --cpu_ddr_clock_bridge/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpu_ddr_clock_bridge_m1_waitrequest AND ((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write));
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line6 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_ddr_clock_bridge_m1_address /= cpu_ddr_clock_bridge_m1_address_last_time))))) = '1' then 
          write(write_line6, now);
          write(write_line6, string'(": "));
          write(write_line6, string'("cpu_ddr_clock_bridge_m1_address did not heed wait!!!"));
          write(output, write_line6.all);
          deallocate (write_line6);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_ddr_clock_bridge_m1_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        cpu_ddr_clock_bridge_m1_byteenable_last_time <= cpu_ddr_clock_bridge_m1_byteenable;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line7 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_ddr_clock_bridge_m1_byteenable /= cpu_ddr_clock_bridge_m1_byteenable_last_time))))) = '1' then 
          write(write_line7, now);
          write(write_line7, string'(": "));
          write(write_line7, string'("cpu_ddr_clock_bridge_m1_byteenable did not heed wait!!!"));
          write(output, write_line7.all);
          deallocate (write_line7);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_ddr_clock_bridge_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_ddr_clock_bridge_m1_read_last_time <= cpu_ddr_clock_bridge_m1_read;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line8 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_ddr_clock_bridge_m1_read) /= std_logic'(cpu_ddr_clock_bridge_m1_read_last_time)))))) = '1' then 
          write(write_line8, now);
          write(write_line8, string'(": "));
          write(write_line8, string'("cpu_ddr_clock_bridge_m1_read did not heed wait!!!"));
          write(output, write_line8.all);
          deallocate (write_line8);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_ddr_clock_bridge_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_ddr_clock_bridge_m1_write_last_time <= cpu_ddr_clock_bridge_m1_write;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line9 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_ddr_clock_bridge_m1_write) /= std_logic'(cpu_ddr_clock_bridge_m1_write_last_time)))))) = '1' then 
          write(write_line9, now);
          write(write_line9, string'(": "));
          write(write_line9, string'("cpu_ddr_clock_bridge_m1_write did not heed wait!!!"));
          write(output, write_line9.all);
          deallocate (write_line9);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_ddr_clock_bridge_m1_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_ddr_clock_bridge_m1_writedata_last_time <= cpu_ddr_clock_bridge_m1_writedata;
      end if;

    end process;

    --cpu_ddr_clock_bridge_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line10 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((cpu_ddr_clock_bridge_m1_writedata /= cpu_ddr_clock_bridge_m1_writedata_last_time)))) AND cpu_ddr_clock_bridge_m1_write)) = '1' then 
          write(write_line10, now);
          write(write_line10, string'(": "));
          write(write_line10, string'("cpu_ddr_clock_bridge_m1_writedata did not heed wait!!!"));
          write(output, write_line10.all);
          deallocate (write_line10);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo read when empty, which is an e_process
    process (clk)
    VARIABLE write_line11 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((empty_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo AND read_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo)) = '1' then 
          write(write_line11, now);
          write(write_line11, string'(": "));
          write(write_line11, string'("cpu_ddr_clock_bridge/m1 negative rdv fifo selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo: read AND empty."));
          write(output, write_line11.all & CR);
          deallocate (write_line11);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo write when full, which is an e_process
    process (clk)
    VARIABLE write_line12 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((full_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo AND write_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo) AND NOT read_selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo)) = '1' then 
          write(write_line12, now);
          write(write_line12, string'(": "));
          write(write_line12, string'("cpu_ddr_clock_bridge/m1 negative rdv fifo selecto_nrdv_cpu_ddr_clock_bridge_m1_1_sdram_s1_fifo: write AND full."));
          write(output, write_line12.all & CR);
          deallocate (write_line12);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cpu_ddr_clock_bridge_bridge_arbitrator is 
end entity cpu_ddr_clock_bridge_bridge_arbitrator;


architecture europa of cpu_ddr_clock_bridge_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity descriptor_memory_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_burstcount : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_chipselect : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_dbs_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_dbs_write_32 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_read : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal d1_descriptor_memory_s1_end_xfer : OUT STD_LOGIC;
                 signal descriptor_memory_s1_address : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal descriptor_memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal descriptor_memory_s1_chipselect : OUT STD_LOGIC;
                 signal descriptor_memory_s1_clken : OUT STD_LOGIC;
                 signal descriptor_memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_memory_s1_reset : OUT STD_LOGIC;
                 signal descriptor_memory_s1_write : OUT STD_LOGIC;
                 signal descriptor_memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1 : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_m1_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC
              );
end entity descriptor_memory_s1_arbitrator;


architecture europa of descriptor_memory_s1_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register_in :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_descriptor_memory_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal descriptor_memory_s1_allgrants :  STD_LOGIC;
                signal descriptor_memory_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal descriptor_memory_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal descriptor_memory_s1_any_continuerequest :  STD_LOGIC;
                signal descriptor_memory_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal descriptor_memory_s1_arb_counter_enable :  STD_LOGIC;
                signal descriptor_memory_s1_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_memory_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_memory_s1_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_memory_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal descriptor_memory_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal descriptor_memory_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal descriptor_memory_s1_begins_xfer :  STD_LOGIC;
                signal descriptor_memory_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_memory_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal descriptor_memory_s1_end_xfer :  STD_LOGIC;
                signal descriptor_memory_s1_firsttransfer :  STD_LOGIC;
                signal descriptor_memory_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal descriptor_memory_s1_in_a_read_cycle :  STD_LOGIC;
                signal descriptor_memory_s1_in_a_write_cycle :  STD_LOGIC;
                signal descriptor_memory_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal descriptor_memory_s1_non_bursting_master_requests :  STD_LOGIC;
                signal descriptor_memory_s1_reg_firsttransfer :  STD_LOGIC;
                signal descriptor_memory_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal descriptor_memory_s1_slavearbiterlockenable :  STD_LOGIC;
                signal descriptor_memory_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal descriptor_memory_s1_unreg_firsttransfer :  STD_LOGIC;
                signal descriptor_memory_s1_waits_for_read :  STD_LOGIC;
                signal descriptor_memory_s1_waits_for_write :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_arbiterlock :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_2 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_3 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_4 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_5 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_6 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_7 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_m1_continuerequest :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register_in :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_saved_grant_descriptor_memory_s1 :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_descriptor_memory_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_descriptor_offset_bridge_m1_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal last_cycle_cpuNios_data_master_granted_slave_descriptor_memory_s1 :  STD_LOGIC;
                signal last_cycle_descriptor_offset_bridge_m1_granted_slave_descriptor_memory_s1 :  STD_LOGIC;
                signal p1_cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register :  STD_LOGIC;
                signal p1_descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register :  STD_LOGIC;
                signal shifted_address_to_descriptor_memory_s1_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal shifted_address_to_descriptor_memory_s1_from_descriptor_offset_bridge_m1 :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_descriptor_memory_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT descriptor_memory_s1_end_xfer;
    end if;

  end process;

  descriptor_memory_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpuNios_data_master_qualified_request_descriptor_memory_s1 OR internal_descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1));
  --assign descriptor_memory_s1_readdata_from_sa = descriptor_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  descriptor_memory_s1_readdata_from_sa <= descriptor_memory_s1_readdata;
  internal_cpuNios_data_master_requests_descriptor_memory_s1 <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 12) & std_logic_vector'("000000000000")) = std_logic_vector'("100000000000010000000000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --registered rdv signal_name registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1 assignment, which is an e_assign
  registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1 <= cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register_in;
  --descriptor_memory_s1_arb_share_counter set values, which is an e_mux
  descriptor_memory_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), std_logic_vector'("00000000000000000000000000000001"))), 4);
  --descriptor_memory_s1_non_bursting_master_requests mux, which is an e_mux
  descriptor_memory_s1_non_bursting_master_requests <= ((internal_cpuNios_data_master_requests_descriptor_memory_s1 OR internal_descriptor_offset_bridge_m1_requests_descriptor_memory_s1) OR internal_cpuNios_data_master_requests_descriptor_memory_s1) OR internal_descriptor_offset_bridge_m1_requests_descriptor_memory_s1;
  --descriptor_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  descriptor_memory_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --descriptor_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  descriptor_memory_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(descriptor_memory_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (descriptor_memory_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(descriptor_memory_s1_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (descriptor_memory_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --descriptor_memory_s1_allgrants all slave grants, which is an e_mux
  descriptor_memory_s1_allgrants <= (((or_reduce(descriptor_memory_s1_grant_vector)) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector));
  --descriptor_memory_s1_end_xfer assignment, which is an e_assign
  descriptor_memory_s1_end_xfer <= NOT ((descriptor_memory_s1_waits_for_read OR descriptor_memory_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_descriptor_memory_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_descriptor_memory_s1 <= descriptor_memory_s1_end_xfer AND (((NOT descriptor_memory_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --descriptor_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  descriptor_memory_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_descriptor_memory_s1 AND descriptor_memory_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_descriptor_memory_s1 AND NOT descriptor_memory_s1_non_bursting_master_requests));
  --descriptor_memory_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_memory_s1_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(descriptor_memory_s1_arb_counter_enable) = '1' then 
        descriptor_memory_s1_arb_share_counter <= descriptor_memory_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --descriptor_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_memory_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(descriptor_memory_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_descriptor_memory_s1)) OR ((end_xfer_arb_share_counter_term_descriptor_memory_s1 AND NOT descriptor_memory_s1_non_bursting_master_requests)))) = '1' then 
        descriptor_memory_s1_slavearbiterlockenable <= or_reduce(descriptor_memory_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpuNios/data_master descriptor_memory/s1 arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= descriptor_memory_s1_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --descriptor_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  descriptor_memory_s1_slavearbiterlockenable2 <= or_reduce(descriptor_memory_s1_arb_share_counter_next_value);
  --cpuNios/data_master descriptor_memory/s1 arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= descriptor_memory_s1_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --descriptor_offset_bridge/m1 descriptor_memory/s1 arbiterlock, which is an e_assign
  descriptor_offset_bridge_m1_arbiterlock <= descriptor_memory_s1_slavearbiterlockenable AND descriptor_offset_bridge_m1_continuerequest;
  --descriptor_offset_bridge/m1 descriptor_memory/s1 arbiterlock2, which is an e_assign
  descriptor_offset_bridge_m1_arbiterlock2 <= descriptor_memory_s1_slavearbiterlockenable2 AND descriptor_offset_bridge_m1_continuerequest;
  --descriptor_offset_bridge/m1 granted descriptor_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_descriptor_offset_bridge_m1_granted_slave_descriptor_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_descriptor_offset_bridge_m1_granted_slave_descriptor_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(descriptor_offset_bridge_m1_saved_grant_descriptor_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_memory_s1_arbitration_holdoff_internal OR NOT internal_descriptor_offset_bridge_m1_requests_descriptor_memory_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_descriptor_offset_bridge_m1_granted_slave_descriptor_memory_s1))))));
    end if;

  end process;

  --descriptor_offset_bridge_m1_continuerequest continued request, which is an e_mux
  descriptor_offset_bridge_m1_continuerequest <= last_cycle_descriptor_offset_bridge_m1_granted_slave_descriptor_memory_s1 AND internal_descriptor_offset_bridge_m1_requests_descriptor_memory_s1;
  --descriptor_memory_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  descriptor_memory_s1_any_continuerequest <= descriptor_offset_bridge_m1_continuerequest OR cpuNios_data_master_continuerequest;
  internal_cpuNios_data_master_qualified_request_descriptor_memory_s1 <= internal_cpuNios_data_master_requests_descriptor_memory_s1 AND NOT (((((cpuNios_data_master_read AND (cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register))) OR (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write))) OR descriptor_offset_bridge_m1_arbiterlock));
  --cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register_in <= ((internal_cpuNios_data_master_granted_descriptor_memory_s1 AND cpuNios_data_master_read) AND NOT descriptor_memory_s1_waits_for_read) AND NOT (cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register);
  --shift register p1 cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register) & A_ToStdLogicVector(cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register_in)));
  --cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register <= p1_cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid cpuNios_data_master_read_data_valid_descriptor_memory_s1, which is an e_mux
  cpuNios_data_master_read_data_valid_descriptor_memory_s1 <= cpuNios_data_master_read_data_valid_descriptor_memory_s1_shift_register;
  --descriptor_memory_s1_writedata mux, which is an e_mux
  descriptor_memory_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_descriptor_memory_s1)) = '1'), cpuNios_data_master_writedata, descriptor_offset_bridge_m1_dbs_write_32);
  --mux descriptor_memory_s1_clken, which is an e_mux
  descriptor_memory_s1_clken <= std_logic'('1');
  internal_descriptor_offset_bridge_m1_requests_descriptor_memory_s1 <= to_std_logic(((Std_Logic_Vector'(descriptor_offset_bridge_m1_address_to_slave(26 DOWNTO 12) & std_logic_vector'("000000000000")) = std_logic_vector'("100000000000010000000000000")))) AND descriptor_offset_bridge_m1_chipselect;
  --cpuNios/data_master granted descriptor_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpuNios_data_master_granted_slave_descriptor_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpuNios_data_master_granted_slave_descriptor_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpuNios_data_master_saved_grant_descriptor_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_memory_s1_arbitration_holdoff_internal OR NOT internal_cpuNios_data_master_requests_descriptor_memory_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpuNios_data_master_granted_slave_descriptor_memory_s1))))));
    end if;

  end process;

  --cpuNios_data_master_continuerequest continued request, which is an e_mux
  cpuNios_data_master_continuerequest <= last_cycle_cpuNios_data_master_granted_slave_descriptor_memory_s1 AND internal_cpuNios_data_master_requests_descriptor_memory_s1;
  internal_descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 <= internal_descriptor_offset_bridge_m1_requests_descriptor_memory_s1 AND NOT (((((NOT(or_reduce(internal_descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1))) AND ((descriptor_offset_bridge_m1_write AND descriptor_offset_bridge_m1_chipselect)))) OR cpuNios_data_master_arbiterlock));
  --descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register_in <= (internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1 AND ((descriptor_offset_bridge_m1_read AND descriptor_offset_bridge_m1_chipselect))) AND NOT descriptor_memory_s1_waits_for_read;
  --shift register p1 descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register) & A_ToStdLogicVector(descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register_in)));
  --descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register <= p1_descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1, which is an e_mux
  descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1 <= descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1_shift_register;
  --allow new arb cycle for descriptor_memory/s1, which is an e_assign
  descriptor_memory_s1_allow_new_arb_cycle <= NOT cpuNios_data_master_arbiterlock AND NOT descriptor_offset_bridge_m1_arbiterlock;
  --descriptor_offset_bridge/m1 assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  descriptor_memory_s1_master_qreq_vector(0) <= internal_descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1;
  --descriptor_offset_bridge/m1 grant descriptor_memory/s1, which is an e_assign
  internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1 <= descriptor_memory_s1_grant_vector(0);
  --descriptor_offset_bridge/m1 saved-grant descriptor_memory/s1, which is an e_assign
  descriptor_offset_bridge_m1_saved_grant_descriptor_memory_s1 <= descriptor_memory_s1_arb_winner(0) AND internal_descriptor_offset_bridge_m1_requests_descriptor_memory_s1;
  --cpuNios/data_master assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  descriptor_memory_s1_master_qreq_vector(1) <= internal_cpuNios_data_master_qualified_request_descriptor_memory_s1;
  --cpuNios/data_master grant descriptor_memory/s1, which is an e_assign
  internal_cpuNios_data_master_granted_descriptor_memory_s1 <= descriptor_memory_s1_grant_vector(1);
  --cpuNios/data_master saved-grant descriptor_memory/s1, which is an e_assign
  cpuNios_data_master_saved_grant_descriptor_memory_s1 <= descriptor_memory_s1_arb_winner(1) AND internal_cpuNios_data_master_requests_descriptor_memory_s1;
  --descriptor_memory/s1 chosen-master double-vector, which is an e_assign
  descriptor_memory_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((descriptor_memory_s1_master_qreq_vector & descriptor_memory_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT descriptor_memory_s1_master_qreq_vector & NOT descriptor_memory_s1_master_qreq_vector))) + (std_logic_vector'("000") & (descriptor_memory_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  descriptor_memory_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((descriptor_memory_s1_allow_new_arb_cycle AND or_reduce(descriptor_memory_s1_grant_vector)))) = '1'), descriptor_memory_s1_grant_vector, descriptor_memory_s1_saved_chosen_master_vector);
  --saved descriptor_memory_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_memory_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(descriptor_memory_s1_allow_new_arb_cycle) = '1' then 
        descriptor_memory_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(descriptor_memory_s1_grant_vector)) = '1'), descriptor_memory_s1_grant_vector, descriptor_memory_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  descriptor_memory_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((descriptor_memory_s1_chosen_master_double_vector(1) OR descriptor_memory_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((descriptor_memory_s1_chosen_master_double_vector(0) OR descriptor_memory_s1_chosen_master_double_vector(2)))));
  --descriptor_memory/s1 chosen master rotated left, which is an e_assign
  descriptor_memory_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(descriptor_memory_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(descriptor_memory_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --descriptor_memory/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_memory_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(descriptor_memory_s1_grant_vector)) = '1' then 
        descriptor_memory_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(descriptor_memory_s1_end_xfer) = '1'), descriptor_memory_s1_chosen_master_rot_left, descriptor_memory_s1_grant_vector);
      end if;
    end if;

  end process;

  --~descriptor_memory_s1_reset assignment, which is an e_assign
  descriptor_memory_s1_reset <= NOT reset_n;
  descriptor_memory_s1_chipselect <= internal_cpuNios_data_master_granted_descriptor_memory_s1 OR internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1;
  --descriptor_memory_s1_firsttransfer first transaction, which is an e_assign
  descriptor_memory_s1_firsttransfer <= A_WE_StdLogic((std_logic'(descriptor_memory_s1_begins_xfer) = '1'), descriptor_memory_s1_unreg_firsttransfer, descriptor_memory_s1_reg_firsttransfer);
  --descriptor_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  descriptor_memory_s1_unreg_firsttransfer <= NOT ((descriptor_memory_s1_slavearbiterlockenable AND descriptor_memory_s1_any_continuerequest));
  --descriptor_memory_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_memory_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(descriptor_memory_s1_begins_xfer) = '1' then 
        descriptor_memory_s1_reg_firsttransfer <= descriptor_memory_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --descriptor_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  descriptor_memory_s1_beginbursttransfer_internal <= descriptor_memory_s1_begins_xfer;
  --descriptor_memory_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  descriptor_memory_s1_arbitration_holdoff_internal <= descriptor_memory_s1_begins_xfer AND descriptor_memory_s1_firsttransfer;
  --descriptor_memory_s1_write assignment, which is an e_mux
  descriptor_memory_s1_write <= ((internal_cpuNios_data_master_granted_descriptor_memory_s1 AND cpuNios_data_master_write)) OR ((internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1 AND ((descriptor_offset_bridge_m1_write AND descriptor_offset_bridge_m1_chipselect))));
  shifted_address_to_descriptor_memory_s1_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --descriptor_memory_s1_address mux, which is an e_mux
  descriptor_memory_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_descriptor_memory_s1)) = '1'), (A_SRL(shifted_address_to_descriptor_memory_s1_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_descriptor_memory_s1_from_descriptor_offset_bridge_m1,std_logic_vector'("00000000000000000000000000000010")))), 10);
  shifted_address_to_descriptor_memory_s1_from_descriptor_offset_bridge_m1 <= A_EXT (Std_Logic_Vector'(A_SRL(descriptor_offset_bridge_m1_address_to_slave,std_logic_vector'("00000000000000000000000000000101")) & descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2) & A_REP(std_logic'('0'), 2)), 27);
  --d1_descriptor_memory_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_descriptor_memory_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_descriptor_memory_s1_end_xfer <= descriptor_memory_s1_end_xfer;
    end if;

  end process;

  --descriptor_memory_s1_waits_for_read in a cycle, which is an e_mux
  descriptor_memory_s1_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_memory_s1_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --descriptor_memory_s1_in_a_read_cycle assignment, which is an e_assign
  descriptor_memory_s1_in_a_read_cycle <= ((internal_cpuNios_data_master_granted_descriptor_memory_s1 AND cpuNios_data_master_read)) OR ((internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1 AND ((descriptor_offset_bridge_m1_read AND descriptor_offset_bridge_m1_chipselect))));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= descriptor_memory_s1_in_a_read_cycle;
  --descriptor_memory_s1_waits_for_write in a cycle, which is an e_mux
  descriptor_memory_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_memory_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --descriptor_memory_s1_in_a_write_cycle assignment, which is an e_assign
  descriptor_memory_s1_in_a_write_cycle <= ((internal_cpuNios_data_master_granted_descriptor_memory_s1 AND cpuNios_data_master_write)) OR ((internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1 AND ((descriptor_offset_bridge_m1_write AND descriptor_offset_bridge_m1_chipselect))));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= descriptor_memory_s1_in_a_write_cycle;
  wait_for_descriptor_memory_s1_counter <= std_logic'('0');
  --descriptor_memory_s1_byteenable byte enable port mux, which is an e_mux
  descriptor_memory_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpuNios_data_master_granted_descriptor_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpuNios_data_master_byteenable)), A_WE_StdLogicVector((std_logic'((internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (internal_descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  (descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_7(3), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_7(2), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_7(1), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_7(0), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_6(3), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_6(2), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_6(1), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_6(0), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_5(3), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_5(2), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_5(1), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_5(0), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_4(3), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_4(2), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_4(1), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_4(0), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_3(3), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_3(2), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_3(1), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_3(0), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_2(3), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_2(2), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_2(1), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_2(0), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_1(3), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_1(2), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_1(1), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_1(0), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_0(3), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_0(2), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_0(1), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_0(0)) <= descriptor_offset_bridge_m1_byteenable;
  internal_descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1 <= A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000000"))), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_0, A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000001"))), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_1, A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000010"))), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_2, A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000011"))), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_3, A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000100"))), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_4, A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000101"))), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_5, A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000110"))), descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_6, descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1_segment_7)))))));
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_descriptor_memory_s1 <= internal_cpuNios_data_master_granted_descriptor_memory_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_descriptor_memory_s1 <= internal_cpuNios_data_master_qualified_request_descriptor_memory_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_descriptor_memory_s1 <= internal_cpuNios_data_master_requests_descriptor_memory_s1;
  --vhdl renameroo for output signals
  descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1 <= internal_descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1;
  --vhdl renameroo for output signals
  descriptor_offset_bridge_m1_granted_descriptor_memory_s1 <= internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1;
  --vhdl renameroo for output signals
  descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 <= internal_descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1;
  --vhdl renameroo for output signals
  descriptor_offset_bridge_m1_requests_descriptor_memory_s1 <= internal_descriptor_offset_bridge_m1_requests_descriptor_memory_s1;
--synthesis translate_off
    --descriptor_memory/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --descriptor_offset_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line13 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_descriptor_offset_bridge_m1_requests_descriptor_memory_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_offset_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line13, now);
          write(write_line13, string'(": "));
          write(write_line13, string'("descriptor_offset_bridge/m1 drove 0 on its 'burstcount' port while accessing slave descriptor_memory/s1"));
          write(output, write_line13.all);
          deallocate (write_line13);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line14 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpuNios_data_master_granted_descriptor_memory_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_descriptor_offset_bridge_m1_granted_descriptor_memory_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line14, now);
          write(write_line14, string'(": "));
          write(write_line14, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line14.all);
          deallocate (write_line14);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line15 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpuNios_data_master_saved_grant_descriptor_memory_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(descriptor_offset_bridge_m1_saved_grant_descriptor_memory_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line15, now);
          write(write_line15, string'(": "));
          write(write_line15, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line15.all);
          deallocate (write_line15);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_sgdma_rx_descriptor_read_to_descriptor_offset_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_sgdma_rx_descriptor_read_to_descriptor_offset_bridge_s1_module;


architecture europa of rdv_fifo_for_sgdma_rx_descriptor_read_to_descriptor_offset_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_sgdma_tx_descriptor_read_to_descriptor_offset_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_sgdma_tx_descriptor_read_to_descriptor_offset_bridge_s1_module;


architecture europa of rdv_fifo_for_sgdma_tx_descriptor_read_to_descriptor_offset_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity descriptor_offset_bridge_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal descriptor_offset_bridge_s1_endofpacket : IN STD_LOGIC;
                 signal descriptor_offset_bridge_s1_readdata : IN STD_LOGIC_VECTOR (255 DOWNTO 0);
                 signal descriptor_offset_bridge_s1_readdatavalid : IN STD_LOGIC;
                 signal descriptor_offset_bridge_s1_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_read_latency_counter : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_read : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_write_write : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_read_latency_counter : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_read : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_write_write : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal d1_descriptor_offset_bridge_s1_end_xfer : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal descriptor_offset_bridge_s1_arbiterlock : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_arbiterlock2 : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_burstcount : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_offset_bridge_s1_chipselect : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_debugaccess : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal descriptor_offset_bridge_s1_read : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (255 DOWNTO 0);
                 signal descriptor_offset_bridge_s1_reset_n : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_write : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (255 DOWNTO 0);
                 signal sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 : OUT STD_LOGIC
              );
end entity descriptor_offset_bridge_s1_arbitrator;


architecture europa of descriptor_offset_bridge_s1_arbitrator is
component rdv_fifo_for_sgdma_rx_descriptor_read_to_descriptor_offset_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_sgdma_rx_descriptor_read_to_descriptor_offset_bridge_s1_module;

component rdv_fifo_for_sgdma_tx_descriptor_read_to_descriptor_offset_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_sgdma_tx_descriptor_read_to_descriptor_offset_bridge_s1_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_allgrants :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_any_continuerequest :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_arb_addend :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_s1_arb_counter_enable :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_arb_share_counter :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_arb_share_set_values :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_arb_winner :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_begins_xfer :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal descriptor_offset_bridge_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_s1_end_xfer :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_firsttransfer :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_grant_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_s1_in_a_read_cycle :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_in_a_write_cycle :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_master_qreq_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_non_bursting_master_requests :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_reg_firsttransfer :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_s1_slavearbiterlockenable :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_unreg_firsttransfer :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_waits_for_read :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_waits_for_write :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_descriptor_offset_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal module_input10 :  STD_LOGIC;
                signal module_input11 :  STD_LOGIC;
                signal module_input12 :  STD_LOGIC;
                signal module_input13 :  STD_LOGIC;
                signal module_input14 :  STD_LOGIC;
                signal module_input9 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_arbiterlock :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_arbiterlock2 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_continuerequest :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_rdv_fifo_empty_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_rdv_fifo_output_from_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_saved_grant_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_arbiterlock :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_arbiterlock2 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_byteenable_descriptor_offset_bridge_s1 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_write_continuerequest :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_saved_grant_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_writedata_replicated :  STD_LOGIC_VECTOR (255 DOWNTO 0);
                signal sgdma_tx_descriptor_read_arbiterlock :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_arbiterlock2 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_continuerequest :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_rdv_fifo_empty_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_rdv_fifo_output_from_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_saved_grant_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_arbiterlock :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_arbiterlock2 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_byteenable_descriptor_offset_bridge_s1 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_write_continuerequest :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_saved_grant_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_writedata_replicated :  STD_LOGIC_VECTOR (255 DOWNTO 0);
                signal shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_rx_descriptor_read :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_rx_descriptor_write :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_tx_descriptor_read :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_tx_descriptor_write :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal wait_for_descriptor_offset_bridge_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT descriptor_offset_bridge_s1_end_xfer;
    end if;

  end process;

  descriptor_offset_bridge_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((((internal_sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 OR internal_sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1));
  --assign descriptor_offset_bridge_s1_readdata_from_sa = descriptor_offset_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  descriptor_offset_bridge_s1_readdata_from_sa <= descriptor_offset_bridge_s1_readdata;
  internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_rx_descriptor_read_address_to_slave(31 DOWNTO 27) & std_logic_vector'("000000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (sgdma_rx_descriptor_read_read))) AND sgdma_rx_descriptor_read_read;
  --assign descriptor_offset_bridge_s1_waitrequest_from_sa = descriptor_offset_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_descriptor_offset_bridge_s1_waitrequest_from_sa <= descriptor_offset_bridge_s1_waitrequest;
  --assign descriptor_offset_bridge_s1_readdatavalid_from_sa = descriptor_offset_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  descriptor_offset_bridge_s1_readdatavalid_from_sa <= descriptor_offset_bridge_s1_readdatavalid;
  --descriptor_offset_bridge_s1_arb_share_counter set values, which is an e_mux
  descriptor_offset_bridge_s1_arb_share_set_values <= std_logic'('1');
  --descriptor_offset_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  descriptor_offset_bridge_s1_non_bursting_master_requests <= ((((((((((((((((((internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 OR internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1) OR internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1) OR internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1) OR internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1) OR internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1) OR internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1) OR internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1) OR internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1) OR internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1;
  --descriptor_offset_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  descriptor_offset_bridge_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --descriptor_offset_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  descriptor_offset_bridge_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(descriptor_offset_bridge_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_offset_bridge_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(descriptor_offset_bridge_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_offset_bridge_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --descriptor_offset_bridge_s1_allgrants all slave grants, which is an e_mux
  descriptor_offset_bridge_s1_allgrants <= (((((((((((((((((((or_reduce(descriptor_offset_bridge_s1_grant_vector)) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector))) OR (or_reduce(descriptor_offset_bridge_s1_grant_vector));
  --descriptor_offset_bridge_s1_end_xfer assignment, which is an e_assign
  descriptor_offset_bridge_s1_end_xfer <= NOT ((descriptor_offset_bridge_s1_waits_for_read OR descriptor_offset_bridge_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_descriptor_offset_bridge_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_descriptor_offset_bridge_s1 <= descriptor_offset_bridge_s1_end_xfer AND (((NOT descriptor_offset_bridge_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --descriptor_offset_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  descriptor_offset_bridge_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_descriptor_offset_bridge_s1 AND descriptor_offset_bridge_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_descriptor_offset_bridge_s1 AND NOT descriptor_offset_bridge_s1_non_bursting_master_requests));
  --descriptor_offset_bridge_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_offset_bridge_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(descriptor_offset_bridge_s1_arb_counter_enable) = '1' then 
        descriptor_offset_bridge_s1_arb_share_counter <= descriptor_offset_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --descriptor_offset_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_offset_bridge_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(descriptor_offset_bridge_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_descriptor_offset_bridge_s1)) OR ((end_xfer_arb_share_counter_term_descriptor_offset_bridge_s1 AND NOT descriptor_offset_bridge_s1_non_bursting_master_requests)))) = '1' then 
        descriptor_offset_bridge_s1_slavearbiterlockenable <= descriptor_offset_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sgdma_rx/descriptor_read descriptor_offset_bridge/s1 arbiterlock, which is an e_assign
  sgdma_rx_descriptor_read_arbiterlock <= descriptor_offset_bridge_s1_slavearbiterlockenable AND sgdma_rx_descriptor_read_continuerequest;
  --descriptor_offset_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  descriptor_offset_bridge_s1_slavearbiterlockenable2 <= descriptor_offset_bridge_s1_arb_share_counter_next_value;
  --sgdma_rx/descriptor_read descriptor_offset_bridge/s1 arbiterlock2, which is an e_assign
  sgdma_rx_descriptor_read_arbiterlock2 <= descriptor_offset_bridge_s1_slavearbiterlockenable2 AND sgdma_rx_descriptor_read_continuerequest;
  --sgdma_rx/descriptor_write descriptor_offset_bridge/s1 arbiterlock, which is an e_assign
  sgdma_rx_descriptor_write_arbiterlock <= descriptor_offset_bridge_s1_slavearbiterlockenable AND sgdma_rx_descriptor_write_continuerequest;
  --sgdma_rx/descriptor_write descriptor_offset_bridge/s1 arbiterlock2, which is an e_assign
  sgdma_rx_descriptor_write_arbiterlock2 <= descriptor_offset_bridge_s1_slavearbiterlockenable2 AND sgdma_rx_descriptor_write_continuerequest;
  --sgdma_rx/descriptor_write granted descriptor_offset_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_rx_descriptor_write_saved_grant_descriptor_offset_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_offset_bridge_s1_arbitration_holdoff_internal OR NOT internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_offset_bridge_s1))))));
    end if;

  end process;

  --sgdma_rx_descriptor_write_continuerequest continued request, which is an e_mux
  sgdma_rx_descriptor_write_continuerequest <= (((last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1)) OR ((last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1))) OR ((last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1));
  --descriptor_offset_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  descriptor_offset_bridge_s1_any_continuerequest <= ((((((((((sgdma_rx_descriptor_write_continuerequest OR sgdma_tx_descriptor_read_continuerequest) OR sgdma_tx_descriptor_write_continuerequest) OR sgdma_rx_descriptor_read_continuerequest) OR sgdma_tx_descriptor_read_continuerequest) OR sgdma_tx_descriptor_write_continuerequest) OR sgdma_rx_descriptor_read_continuerequest) OR sgdma_rx_descriptor_write_continuerequest) OR sgdma_tx_descriptor_write_continuerequest) OR sgdma_rx_descriptor_read_continuerequest) OR sgdma_rx_descriptor_write_continuerequest) OR sgdma_tx_descriptor_read_continuerequest;
  --sgdma_tx/descriptor_read descriptor_offset_bridge/s1 arbiterlock, which is an e_assign
  sgdma_tx_descriptor_read_arbiterlock <= descriptor_offset_bridge_s1_slavearbiterlockenable AND sgdma_tx_descriptor_read_continuerequest;
  --sgdma_tx/descriptor_read descriptor_offset_bridge/s1 arbiterlock2, which is an e_assign
  sgdma_tx_descriptor_read_arbiterlock2 <= descriptor_offset_bridge_s1_slavearbiterlockenable2 AND sgdma_tx_descriptor_read_continuerequest;
  --sgdma_tx/descriptor_read granted descriptor_offset_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_tx_descriptor_read_saved_grant_descriptor_offset_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_offset_bridge_s1_arbitration_holdoff_internal OR NOT internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_offset_bridge_s1))))));
    end if;

  end process;

  --sgdma_tx_descriptor_read_continuerequest continued request, which is an e_mux
  sgdma_tx_descriptor_read_continuerequest <= (((last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1)) OR ((last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1))) OR ((last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1));
  --sgdma_tx/descriptor_write descriptor_offset_bridge/s1 arbiterlock, which is an e_assign
  sgdma_tx_descriptor_write_arbiterlock <= descriptor_offset_bridge_s1_slavearbiterlockenable AND sgdma_tx_descriptor_write_continuerequest;
  --sgdma_tx/descriptor_write descriptor_offset_bridge/s1 arbiterlock2, which is an e_assign
  sgdma_tx_descriptor_write_arbiterlock2 <= descriptor_offset_bridge_s1_slavearbiterlockenable2 AND sgdma_tx_descriptor_write_continuerequest;
  --sgdma_tx/descriptor_write granted descriptor_offset_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_tx_descriptor_write_saved_grant_descriptor_offset_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_offset_bridge_s1_arbitration_holdoff_internal OR NOT internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_offset_bridge_s1))))));
    end if;

  end process;

  --sgdma_tx_descriptor_write_continuerequest continued request, which is an e_mux
  sgdma_tx_descriptor_write_continuerequest <= (((last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1)) OR ((last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1))) OR ((last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1));
  internal_sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 <= internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 AND NOT ((((((sgdma_rx_descriptor_read_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_rx_descriptor_read_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_rx_descriptor_read_latency_counter)))))))))) OR sgdma_rx_descriptor_write_arbiterlock) OR sgdma_tx_descriptor_read_arbiterlock) OR sgdma_tx_descriptor_write_arbiterlock));
  --unique name for descriptor_offset_bridge_s1_move_on_to_next_transaction, which is an e_assign
  descriptor_offset_bridge_s1_move_on_to_next_transaction <= descriptor_offset_bridge_s1_readdatavalid_from_sa;
  --rdv_fifo_for_sgdma_rx_descriptor_read_to_descriptor_offset_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_sgdma_rx_descriptor_read_to_descriptor_offset_bridge_s1 : rdv_fifo_for_sgdma_rx_descriptor_read_to_descriptor_offset_bridge_s1_module
    port map(
      data_out => sgdma_rx_descriptor_read_rdv_fifo_output_from_descriptor_offset_bridge_s1,
      empty => open,
      fifo_contains_ones_n => sgdma_rx_descriptor_read_rdv_fifo_empty_descriptor_offset_bridge_s1,
      full => open,
      clear_fifo => module_input9,
      clk => clk,
      data_in => internal_sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1,
      read => descriptor_offset_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input10,
      write => module_input11
    );

  module_input9 <= std_logic'('0');
  module_input10 <= std_logic'('0');
  module_input11 <= in_a_read_cycle AND NOT descriptor_offset_bridge_s1_waits_for_read;

  sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register <= NOT sgdma_rx_descriptor_read_rdv_fifo_empty_descriptor_offset_bridge_s1;
  --local readdatavalid sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1, which is an e_mux
  sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 <= ((descriptor_offset_bridge_s1_readdatavalid_from_sa AND sgdma_rx_descriptor_read_rdv_fifo_output_from_descriptor_offset_bridge_s1)) AND NOT sgdma_rx_descriptor_read_rdv_fifo_empty_descriptor_offset_bridge_s1;
  --assign descriptor_offset_bridge_s1_endofpacket_from_sa = descriptor_offset_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  descriptor_offset_bridge_s1_endofpacket_from_sa <= descriptor_offset_bridge_s1_endofpacket;
  internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_rx_descriptor_write_address_to_slave(31 DOWNTO 27) & std_logic_vector'("000000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (sgdma_rx_descriptor_write_write))) AND sgdma_rx_descriptor_write_write;
  --sgdma_rx/descriptor_read granted descriptor_offset_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_rx_descriptor_read_saved_grant_descriptor_offset_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_offset_bridge_s1_arbitration_holdoff_internal OR NOT internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_offset_bridge_s1))))));
    end if;

  end process;

  --sgdma_rx_descriptor_read_continuerequest continued request, which is an e_mux
  sgdma_rx_descriptor_read_continuerequest <= (((last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1)) OR ((last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1))) OR ((last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_offset_bridge_s1 AND internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1));
  internal_sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 <= internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 AND NOT (((sgdma_rx_descriptor_read_arbiterlock OR sgdma_tx_descriptor_read_arbiterlock) OR sgdma_tx_descriptor_write_arbiterlock));
  --replicate narrow data for wide slave
  sgdma_rx_descriptor_write_writedata_replicated <= sgdma_rx_descriptor_write_writedata & sgdma_rx_descriptor_write_writedata & sgdma_rx_descriptor_write_writedata & sgdma_rx_descriptor_write_writedata & sgdma_rx_descriptor_write_writedata & sgdma_rx_descriptor_write_writedata & sgdma_rx_descriptor_write_writedata & sgdma_rx_descriptor_write_writedata;
  --descriptor_offset_bridge_s1_writedata mux, which is an e_mux
  descriptor_offset_bridge_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1)) = '1'), sgdma_rx_descriptor_write_writedata_replicated, sgdma_tx_descriptor_write_writedata_replicated);
  internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_tx_descriptor_read_address_to_slave(31 DOWNTO 27) & std_logic_vector'("000000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (sgdma_tx_descriptor_read_read))) AND sgdma_tx_descriptor_read_read;
  internal_sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 <= internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 AND NOT ((((((sgdma_tx_descriptor_read_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_tx_descriptor_read_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_tx_descriptor_read_latency_counter)))))))))) OR sgdma_rx_descriptor_read_arbiterlock) OR sgdma_rx_descriptor_write_arbiterlock) OR sgdma_tx_descriptor_write_arbiterlock));
  --rdv_fifo_for_sgdma_tx_descriptor_read_to_descriptor_offset_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_sgdma_tx_descriptor_read_to_descriptor_offset_bridge_s1 : rdv_fifo_for_sgdma_tx_descriptor_read_to_descriptor_offset_bridge_s1_module
    port map(
      data_out => sgdma_tx_descriptor_read_rdv_fifo_output_from_descriptor_offset_bridge_s1,
      empty => open,
      fifo_contains_ones_n => sgdma_tx_descriptor_read_rdv_fifo_empty_descriptor_offset_bridge_s1,
      full => open,
      clear_fifo => module_input12,
      clk => clk,
      data_in => internal_sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1,
      read => descriptor_offset_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input13,
      write => module_input14
    );

  module_input12 <= std_logic'('0');
  module_input13 <= std_logic'('0');
  module_input14 <= in_a_read_cycle AND NOT descriptor_offset_bridge_s1_waits_for_read;

  sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register <= NOT sgdma_tx_descriptor_read_rdv_fifo_empty_descriptor_offset_bridge_s1;
  --local readdatavalid sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1, which is an e_mux
  sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 <= ((descriptor_offset_bridge_s1_readdatavalid_from_sa AND sgdma_tx_descriptor_read_rdv_fifo_output_from_descriptor_offset_bridge_s1)) AND NOT sgdma_tx_descriptor_read_rdv_fifo_empty_descriptor_offset_bridge_s1;
  internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_tx_descriptor_write_address_to_slave(31 DOWNTO 27) & std_logic_vector'("000000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (sgdma_tx_descriptor_write_write))) AND sgdma_tx_descriptor_write_write;
  internal_sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 <= internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 AND NOT (((sgdma_rx_descriptor_read_arbiterlock OR sgdma_rx_descriptor_write_arbiterlock) OR sgdma_tx_descriptor_read_arbiterlock));
  --replicate narrow data for wide slave
  sgdma_tx_descriptor_write_writedata_replicated <= sgdma_tx_descriptor_write_writedata & sgdma_tx_descriptor_write_writedata & sgdma_tx_descriptor_write_writedata & sgdma_tx_descriptor_write_writedata & sgdma_tx_descriptor_write_writedata & sgdma_tx_descriptor_write_writedata & sgdma_tx_descriptor_write_writedata & sgdma_tx_descriptor_write_writedata;
  --allow new arb cycle for descriptor_offset_bridge/s1, which is an e_assign
  descriptor_offset_bridge_s1_allow_new_arb_cycle <= ((NOT sgdma_rx_descriptor_read_arbiterlock AND NOT sgdma_rx_descriptor_write_arbiterlock) AND NOT sgdma_tx_descriptor_read_arbiterlock) AND NOT sgdma_tx_descriptor_write_arbiterlock;
  --sgdma_tx/descriptor_write assignment into master qualified-requests vector for descriptor_offset_bridge/s1, which is an e_assign
  descriptor_offset_bridge_s1_master_qreq_vector(0) <= internal_sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1;
  --sgdma_tx/descriptor_write grant descriptor_offset_bridge/s1, which is an e_assign
  internal_sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 <= descriptor_offset_bridge_s1_grant_vector(0);
  --sgdma_tx/descriptor_write saved-grant descriptor_offset_bridge/s1, which is an e_assign
  sgdma_tx_descriptor_write_saved_grant_descriptor_offset_bridge_s1 <= descriptor_offset_bridge_s1_arb_winner(0) AND internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1;
  --sgdma_tx/descriptor_read assignment into master qualified-requests vector for descriptor_offset_bridge/s1, which is an e_assign
  descriptor_offset_bridge_s1_master_qreq_vector(1) <= internal_sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1;
  --sgdma_tx/descriptor_read grant descriptor_offset_bridge/s1, which is an e_assign
  internal_sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 <= descriptor_offset_bridge_s1_grant_vector(1);
  --sgdma_tx/descriptor_read saved-grant descriptor_offset_bridge/s1, which is an e_assign
  sgdma_tx_descriptor_read_saved_grant_descriptor_offset_bridge_s1 <= descriptor_offset_bridge_s1_arb_winner(1) AND internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1;
  --sgdma_rx/descriptor_write assignment into master qualified-requests vector for descriptor_offset_bridge/s1, which is an e_assign
  descriptor_offset_bridge_s1_master_qreq_vector(2) <= internal_sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1;
  --sgdma_rx/descriptor_write grant descriptor_offset_bridge/s1, which is an e_assign
  internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 <= descriptor_offset_bridge_s1_grant_vector(2);
  --sgdma_rx/descriptor_write saved-grant descriptor_offset_bridge/s1, which is an e_assign
  sgdma_rx_descriptor_write_saved_grant_descriptor_offset_bridge_s1 <= descriptor_offset_bridge_s1_arb_winner(2) AND internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1;
  --sgdma_rx/descriptor_read assignment into master qualified-requests vector for descriptor_offset_bridge/s1, which is an e_assign
  descriptor_offset_bridge_s1_master_qreq_vector(3) <= internal_sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1;
  --sgdma_rx/descriptor_read grant descriptor_offset_bridge/s1, which is an e_assign
  internal_sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 <= descriptor_offset_bridge_s1_grant_vector(3);
  --sgdma_rx/descriptor_read saved-grant descriptor_offset_bridge/s1, which is an e_assign
  sgdma_rx_descriptor_read_saved_grant_descriptor_offset_bridge_s1 <= descriptor_offset_bridge_s1_arb_winner(3) AND internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1;
  --descriptor_offset_bridge/s1 chosen-master double-vector, which is an e_assign
  descriptor_offset_bridge_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((descriptor_offset_bridge_s1_master_qreq_vector & descriptor_offset_bridge_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT descriptor_offset_bridge_s1_master_qreq_vector & NOT descriptor_offset_bridge_s1_master_qreq_vector))) + (std_logic_vector'("00000") & (descriptor_offset_bridge_s1_arb_addend))))), 8);
  --stable onehot encoding of arb winner
  descriptor_offset_bridge_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((descriptor_offset_bridge_s1_allow_new_arb_cycle AND or_reduce(descriptor_offset_bridge_s1_grant_vector)))) = '1'), descriptor_offset_bridge_s1_grant_vector, descriptor_offset_bridge_s1_saved_chosen_master_vector);
  --saved descriptor_offset_bridge_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_offset_bridge_s1_saved_chosen_master_vector <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(descriptor_offset_bridge_s1_allow_new_arb_cycle) = '1' then 
        descriptor_offset_bridge_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(descriptor_offset_bridge_s1_grant_vector)) = '1'), descriptor_offset_bridge_s1_grant_vector, descriptor_offset_bridge_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  descriptor_offset_bridge_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((descriptor_offset_bridge_s1_chosen_master_double_vector(3) OR descriptor_offset_bridge_s1_chosen_master_double_vector(7)))) & A_ToStdLogicVector(((descriptor_offset_bridge_s1_chosen_master_double_vector(2) OR descriptor_offset_bridge_s1_chosen_master_double_vector(6)))) & A_ToStdLogicVector(((descriptor_offset_bridge_s1_chosen_master_double_vector(1) OR descriptor_offset_bridge_s1_chosen_master_double_vector(5)))) & A_ToStdLogicVector(((descriptor_offset_bridge_s1_chosen_master_double_vector(0) OR descriptor_offset_bridge_s1_chosen_master_double_vector(4)))));
  --descriptor_offset_bridge/s1 chosen master rotated left, which is an e_assign
  descriptor_offset_bridge_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(descriptor_offset_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("0000")), (std_logic_vector'("0000000000000000000000000000") & ((A_SLL(descriptor_offset_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 4);
  --descriptor_offset_bridge/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_offset_bridge_s1_arb_addend <= std_logic_vector'("0001");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(descriptor_offset_bridge_s1_grant_vector)) = '1' then 
        descriptor_offset_bridge_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(descriptor_offset_bridge_s1_end_xfer) = '1'), descriptor_offset_bridge_s1_chosen_master_rot_left, descriptor_offset_bridge_s1_grant_vector);
      end if;
    end if;

  end process;

  --descriptor_offset_bridge_s1_reset_n assignment, which is an e_assign
  descriptor_offset_bridge_s1_reset_n <= reset_n;
  descriptor_offset_bridge_s1_chipselect <= ((internal_sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 OR internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1) OR internal_sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1;
  --descriptor_offset_bridge_s1_firsttransfer first transaction, which is an e_assign
  descriptor_offset_bridge_s1_firsttransfer <= A_WE_StdLogic((std_logic'(descriptor_offset_bridge_s1_begins_xfer) = '1'), descriptor_offset_bridge_s1_unreg_firsttransfer, descriptor_offset_bridge_s1_reg_firsttransfer);
  --descriptor_offset_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  descriptor_offset_bridge_s1_unreg_firsttransfer <= NOT ((descriptor_offset_bridge_s1_slavearbiterlockenable AND descriptor_offset_bridge_s1_any_continuerequest));
  --descriptor_offset_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_offset_bridge_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(descriptor_offset_bridge_s1_begins_xfer) = '1' then 
        descriptor_offset_bridge_s1_reg_firsttransfer <= descriptor_offset_bridge_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --descriptor_offset_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  descriptor_offset_bridge_s1_beginbursttransfer_internal <= descriptor_offset_bridge_s1_begins_xfer;
  --descriptor_offset_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  descriptor_offset_bridge_s1_arbitration_holdoff_internal <= descriptor_offset_bridge_s1_begins_xfer AND descriptor_offset_bridge_s1_firsttransfer;
  --descriptor_offset_bridge_s1_read assignment, which is an e_mux
  descriptor_offset_bridge_s1_read <= ((internal_sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 AND sgdma_rx_descriptor_read_read)) OR ((internal_sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 AND sgdma_tx_descriptor_read_read));
  --descriptor_offset_bridge_s1_write assignment, which is an e_mux
  descriptor_offset_bridge_s1_write <= ((internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 AND sgdma_rx_descriptor_write_write)) OR ((internal_sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 AND sgdma_tx_descriptor_write_write));
  shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_rx_descriptor_read <= sgdma_rx_descriptor_read_address_to_slave;
  --descriptor_offset_bridge_s1_address mux, which is an e_mux
  descriptor_offset_bridge_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1)) = '1'), (A_SRL(shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_rx_descriptor_read,std_logic_vector'("00000000000000000000000000000101"))), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1)) = '1'), (A_SRL(shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_rx_descriptor_write,std_logic_vector'("00000000000000000000000000000101"))), A_WE_StdLogicVector((std_logic'((internal_sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1)) = '1'), (A_SRL(shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_tx_descriptor_read,std_logic_vector'("00000000000000000000000000000101"))), (A_SRL(shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_tx_descriptor_write,std_logic_vector'("00000000000000000000000000000101")))))), 22);
  shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_rx_descriptor_write <= sgdma_rx_descriptor_write_address_to_slave;
  shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_tx_descriptor_read <= sgdma_tx_descriptor_read_address_to_slave;
  shifted_address_to_descriptor_offset_bridge_s1_from_sgdma_tx_descriptor_write <= sgdma_tx_descriptor_write_address_to_slave;
  --slaveid descriptor_offset_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  descriptor_offset_bridge_s1_nativeaddress <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1)) = '1'), (A_SRL(sgdma_rx_descriptor_read_address_to_slave,std_logic_vector'("00000000000000000000000000000010"))), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1)) = '1'), (A_SRL(sgdma_rx_descriptor_write_address_to_slave,std_logic_vector'("00000000000000000000000000000010"))), A_WE_StdLogicVector((std_logic'((internal_sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1)) = '1'), (A_SRL(sgdma_tx_descriptor_read_address_to_slave,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(sgdma_tx_descriptor_write_address_to_slave,std_logic_vector'("00000000000000000000000000000010")))))), 22);
  --d1_descriptor_offset_bridge_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_descriptor_offset_bridge_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_descriptor_offset_bridge_s1_end_xfer <= descriptor_offset_bridge_s1_end_xfer;
    end if;

  end process;

  --descriptor_offset_bridge_s1_waits_for_read in a cycle, which is an e_mux
  descriptor_offset_bridge_s1_waits_for_read <= descriptor_offset_bridge_s1_in_a_read_cycle AND internal_descriptor_offset_bridge_s1_waitrequest_from_sa;
  --descriptor_offset_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  descriptor_offset_bridge_s1_in_a_read_cycle <= ((internal_sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 AND sgdma_rx_descriptor_read_read)) OR ((internal_sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 AND sgdma_tx_descriptor_read_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= descriptor_offset_bridge_s1_in_a_read_cycle;
  --descriptor_offset_bridge_s1_waits_for_write in a cycle, which is an e_mux
  descriptor_offset_bridge_s1_waits_for_write <= descriptor_offset_bridge_s1_in_a_write_cycle AND internal_descriptor_offset_bridge_s1_waitrequest_from_sa;
  --descriptor_offset_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  descriptor_offset_bridge_s1_in_a_write_cycle <= ((internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 AND sgdma_rx_descriptor_write_write)) OR ((internal_sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 AND sgdma_tx_descriptor_write_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= descriptor_offset_bridge_s1_in_a_write_cycle;
  wait_for_descriptor_offset_bridge_s1_counter <= std_logic'('0');
  --descriptor_offset_bridge_s1_byteenable byte enable port mux, which is an e_mux
  descriptor_offset_bridge_s1_byteenable <= A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1)) = '1'), sgdma_rx_descriptor_write_byteenable_descriptor_offset_bridge_s1, A_WE_StdLogicVector((std_logic'((internal_sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1)) = '1'), sgdma_tx_descriptor_write_byteenable_descriptor_offset_bridge_s1, -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --byte_enable_mux for sgdma_rx/descriptor_write and descriptor_offset_bridge/s1, which is an e_mux
  sgdma_rx_descriptor_write_byteenable_descriptor_offset_bridge_s1 <= A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_rx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000") & (A_REP(std_logic'('1'), 4))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_rx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000001"))), (std_logic_vector'("000000000000000000000000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("0000")))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_rx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000010"))), (std_logic_vector'("00000000000000000000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("00000000")))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_rx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000011"))), (std_logic_vector'("0000000000000000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("000000000000")))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_rx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000100"))), (std_logic_vector'("000000000000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("0000000000000000")))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_rx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000101"))), (std_logic_vector'("00000000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("00000000000000000000")))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_rx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000110"))), (std_logic_vector'("0000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("000000000000000000000000")))), (A_REP(std_logic'('1'), 4) & std_logic_vector'("0000000000000000000000000000")))))))));
  --byte_enable_mux for sgdma_tx/descriptor_write and descriptor_offset_bridge/s1, which is an e_mux
  sgdma_tx_descriptor_write_byteenable_descriptor_offset_bridge_s1 <= A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000") & (A_REP(std_logic'('1'), 4))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000001"))), (std_logic_vector'("000000000000000000000000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("0000")))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000010"))), (std_logic_vector'("00000000000000000000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("00000000")))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000011"))), (std_logic_vector'("0000000000000000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("000000000000")))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000100"))), (std_logic_vector'("000000000000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("0000000000000000")))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000101"))), (std_logic_vector'("00000000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("00000000000000000000")))), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_descriptor_write_address_to_slave(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000110"))), (std_logic_vector'("0000") & ((A_REP(std_logic'('1'), 4) & std_logic_vector'("000000000000000000000000")))), (A_REP(std_logic'('1'), 4) & std_logic_vector'("0000000000000000000000000000")))))))));
  --burstcount mux, which is an e_mux
  descriptor_offset_bridge_s1_burstcount <= std_logic'('1');
  --descriptor_offset_bridge/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  descriptor_offset_bridge_s1_arbiterlock <= A_WE_StdLogic((std_logic'((sgdma_rx_descriptor_read_arbiterlock)) = '1'), sgdma_rx_descriptor_read_arbiterlock, A_WE_StdLogic((std_logic'((sgdma_rx_descriptor_write_arbiterlock)) = '1'), sgdma_rx_descriptor_write_arbiterlock, A_WE_StdLogic((std_logic'((sgdma_tx_descriptor_read_arbiterlock)) = '1'), sgdma_tx_descriptor_read_arbiterlock, sgdma_tx_descriptor_write_arbiterlock)));
  --descriptor_offset_bridge/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  descriptor_offset_bridge_s1_arbiterlock2 <= A_WE_StdLogic((std_logic'((sgdma_rx_descriptor_read_arbiterlock2)) = '1'), sgdma_rx_descriptor_read_arbiterlock2, A_WE_StdLogic((std_logic'((sgdma_rx_descriptor_write_arbiterlock2)) = '1'), sgdma_rx_descriptor_write_arbiterlock2, A_WE_StdLogic((std_logic'((sgdma_tx_descriptor_read_arbiterlock2)) = '1'), sgdma_tx_descriptor_read_arbiterlock2, sgdma_tx_descriptor_write_arbiterlock2)));
  --debugaccess mux, which is an e_mux
  descriptor_offset_bridge_s1_debugaccess <= std_logic'('0');
  --vhdl renameroo for output signals
  descriptor_offset_bridge_s1_waitrequest_from_sa <= internal_descriptor_offset_bridge_s1_waitrequest_from_sa;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 <= internal_sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 <= internal_sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 <= internal_sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 <= internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 <= internal_sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 <= internal_sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 <= internal_sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 <= internal_sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 <= internal_sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 <= internal_sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 <= internal_sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 <= internal_sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1;
--synthesis translate_off
    --descriptor_offset_bridge/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line16 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("0000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line16, now);
          write(write_line16, string'(": "));
          write(write_line16, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line16.all);
          deallocate (write_line16);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line17 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("0000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(sgdma_rx_descriptor_read_saved_grant_descriptor_offset_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(sgdma_rx_descriptor_write_saved_grant_descriptor_offset_bridge_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(sgdma_tx_descriptor_read_saved_grant_descriptor_offset_bridge_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(sgdma_tx_descriptor_write_saved_grant_descriptor_offset_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line17, now);
          write(write_line17, string'(": "));
          write(write_line17, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line17.all);
          deallocate (write_line17);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity descriptor_offset_bridge_m1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                 signal descriptor_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_address : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_burstcount : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1 : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_chipselect : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_granted_descriptor_memory_s1 : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_read : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_requests_descriptor_memory_s1 : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_write : IN STD_LOGIC;
                 signal descriptor_offset_bridge_m1_writedata : IN STD_LOGIC_VECTOR (255 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal descriptor_offset_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_dbs_address : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_dbs_write_32 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_latency_counter : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (255 DOWNTO 0);
                 signal descriptor_offset_bridge_m1_readdatavalid : OUT STD_LOGIC;
                 signal descriptor_offset_bridge_m1_waitrequest : OUT STD_LOGIC
              );
end entity descriptor_offset_bridge_m1_arbitrator;


architecture europa of descriptor_offset_bridge_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_32_reg_segment_0 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_latent_32_reg_segment_1 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_latent_32_reg_segment_2 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_latent_32_reg_segment_3 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_latent_32_reg_segment_4 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_latent_32_reg_segment_5 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_latent_32_reg_segment_6 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_address_last_time :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal descriptor_offset_bridge_m1_burstcount_last_time :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_byteenable_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal descriptor_offset_bridge_m1_chipselect_last_time :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_dbs_increment :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_offset_bridge_m1_dbs_rdv_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_offset_bridge_m1_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_offset_bridge_m1_is_granted_some_slave :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_offset_bridge_m1_read_but_no_slave_selected :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_read_last_time :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_run :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_write_last_time :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_writedata_last_time :  STD_LOGIC_VECTOR (255 DOWNTO 0);
                signal internal_descriptor_offset_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal internal_descriptor_offset_bridge_m1_dbs_address :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal internal_descriptor_offset_bridge_m1_latency_counter :  STD_LOGIC;
                signal internal_descriptor_offset_bridge_m1_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p1_dbs_latent_32_reg_segment_0 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_dbs_latent_32_reg_segment_1 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_dbs_latent_32_reg_segment_2 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_dbs_latent_32_reg_segment_3 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_dbs_latent_32_reg_segment_4 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_dbs_latent_32_reg_segment_5 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_dbs_latent_32_reg_segment_6 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_descriptor_offset_bridge_m1_latency_counter :  STD_LOGIC;
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_descriptor_offset_bridge_m1_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 OR (((((((descriptor_offset_bridge_m1_write AND descriptor_offset_bridge_m1_chipselect)) AND NOT(or_reduce(descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1))) AND internal_descriptor_offset_bridge_m1_dbs_address(4)) AND internal_descriptor_offset_bridge_m1_dbs_address(3)) AND internal_descriptor_offset_bridge_m1_dbs_address(2)))) OR NOT descriptor_offset_bridge_m1_requests_descriptor_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((descriptor_offset_bridge_m1_granted_descriptor_memory_s1 OR NOT descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 OR NOT ((descriptor_offset_bridge_m1_read AND descriptor_offset_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((internal_descriptor_offset_bridge_m1_dbs_address(4) AND internal_descriptor_offset_bridge_m1_dbs_address(3)) AND internal_descriptor_offset_bridge_m1_dbs_address(2))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((descriptor_offset_bridge_m1_read AND descriptor_offset_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 OR NOT ((descriptor_offset_bridge_m1_write AND descriptor_offset_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((internal_descriptor_offset_bridge_m1_dbs_address(4) AND internal_descriptor_offset_bridge_m1_dbs_address(3)) AND internal_descriptor_offset_bridge_m1_dbs_address(2))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((descriptor_offset_bridge_m1_write AND descriptor_offset_bridge_m1_chipselect)))))))))));
  --cascaded wait assignment, which is an e_assign
  descriptor_offset_bridge_m1_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_descriptor_offset_bridge_m1_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("100000000000010") & descriptor_offset_bridge_m1_address(11 DOWNTO 0));
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic((((((((NOT std_logic_vector'("00000000000000000000000000000000")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_offset_bridge_m1_requests_descriptor_memory_s1)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((descriptor_offset_bridge_m1_write AND descriptor_offset_bridge_m1_chipselect)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT(or_reduce(descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1))))))) OR ((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((descriptor_offset_bridge_m1_granted_descriptor_memory_s1 AND ((descriptor_offset_bridge_m1_read AND descriptor_offset_bridge_m1_chipselect)))))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")))) OR ((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((descriptor_offset_bridge_m1_granted_descriptor_memory_s1 AND ((descriptor_offset_bridge_m1_write AND descriptor_offset_bridge_m1_chipselect)))))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")))));
  --descriptor_offset_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_offset_bridge_m1_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      descriptor_offset_bridge_m1_read_but_no_slave_selected <= (((descriptor_offset_bridge_m1_read AND descriptor_offset_bridge_m1_chipselect)) AND descriptor_offset_bridge_m1_run) AND NOT descriptor_offset_bridge_m1_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  descriptor_offset_bridge_m1_is_granted_some_slave <= descriptor_offset_bridge_m1_granted_descriptor_memory_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_descriptor_offset_bridge_m1_readdatavalid <= descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1 AND dbs_rdv_counter_overflow;
  --latent slave read data valid which is not flushed, which is an e_mux
  descriptor_offset_bridge_m1_readdatavalid <= descriptor_offset_bridge_m1_read_but_no_slave_selected OR pre_flush_descriptor_offset_bridge_m1_readdatavalid;
  --input to latent dbs-32 stored 0, which is an e_mux
  p1_dbs_latent_32_reg_segment_0 <= descriptor_memory_s1_readdata_from_sa;
  --dbs register for latent dbs-32 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_32_reg_segment_0 <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & ((descriptor_offset_bridge_m1_dbs_rdv_counter(4 DOWNTO 2)))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_32_reg_segment_0 <= p1_dbs_latent_32_reg_segment_0;
      end if;
    end if;

  end process;

  --input to latent dbs-32 stored 1, which is an e_mux
  p1_dbs_latent_32_reg_segment_1 <= descriptor_memory_s1_readdata_from_sa;
  --dbs register for latent dbs-32 segment 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_32_reg_segment_1 <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & ((descriptor_offset_bridge_m1_dbs_rdv_counter(4 DOWNTO 2)))) = std_logic_vector'("00000000000000000000000000000001")))))) = '1' then 
        dbs_latent_32_reg_segment_1 <= p1_dbs_latent_32_reg_segment_1;
      end if;
    end if;

  end process;

  --input to latent dbs-32 stored 2, which is an e_mux
  p1_dbs_latent_32_reg_segment_2 <= descriptor_memory_s1_readdata_from_sa;
  --dbs register for latent dbs-32 segment 2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_32_reg_segment_2 <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & ((descriptor_offset_bridge_m1_dbs_rdv_counter(4 DOWNTO 2)))) = std_logic_vector'("00000000000000000000000000000010")))))) = '1' then 
        dbs_latent_32_reg_segment_2 <= p1_dbs_latent_32_reg_segment_2;
      end if;
    end if;

  end process;

  --input to latent dbs-32 stored 3, which is an e_mux
  p1_dbs_latent_32_reg_segment_3 <= descriptor_memory_s1_readdata_from_sa;
  --dbs register for latent dbs-32 segment 3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_32_reg_segment_3 <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & ((descriptor_offset_bridge_m1_dbs_rdv_counter(4 DOWNTO 2)))) = std_logic_vector'("00000000000000000000000000000011")))))) = '1' then 
        dbs_latent_32_reg_segment_3 <= p1_dbs_latent_32_reg_segment_3;
      end if;
    end if;

  end process;

  --input to latent dbs-32 stored 4, which is an e_mux
  p1_dbs_latent_32_reg_segment_4 <= descriptor_memory_s1_readdata_from_sa;
  --dbs register for latent dbs-32 segment 4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_32_reg_segment_4 <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & ((descriptor_offset_bridge_m1_dbs_rdv_counter(4 DOWNTO 2)))) = std_logic_vector'("00000000000000000000000000000100")))))) = '1' then 
        dbs_latent_32_reg_segment_4 <= p1_dbs_latent_32_reg_segment_4;
      end if;
    end if;

  end process;

  --input to latent dbs-32 stored 5, which is an e_mux
  p1_dbs_latent_32_reg_segment_5 <= descriptor_memory_s1_readdata_from_sa;
  --dbs register for latent dbs-32 segment 5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_32_reg_segment_5 <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & ((descriptor_offset_bridge_m1_dbs_rdv_counter(4 DOWNTO 2)))) = std_logic_vector'("00000000000000000000000000000101")))))) = '1' then 
        dbs_latent_32_reg_segment_5 <= p1_dbs_latent_32_reg_segment_5;
      end if;
    end if;

  end process;

  --input to latent dbs-32 stored 6, which is an e_mux
  p1_dbs_latent_32_reg_segment_6 <= descriptor_memory_s1_readdata_from_sa;
  --dbs register for latent dbs-32 segment 6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_32_reg_segment_6 <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("00000000000000000000000000000") & ((descriptor_offset_bridge_m1_dbs_rdv_counter(4 DOWNTO 2)))) = std_logic_vector'("00000000000000000000000000000110")))))) = '1' then 
        dbs_latent_32_reg_segment_6 <= p1_dbs_latent_32_reg_segment_6;
      end if;
    end if;

  end process;

  --descriptor_offset_bridge/m1 readdata mux, which is an e_mux
  descriptor_offset_bridge_m1_readdata <= Std_Logic_Vector'(descriptor_memory_s1_readdata_from_sa(31 DOWNTO 0) & dbs_latent_32_reg_segment_6 & dbs_latent_32_reg_segment_5 & dbs_latent_32_reg_segment_4 & dbs_latent_32_reg_segment_3 & dbs_latent_32_reg_segment_2 & dbs_latent_32_reg_segment_1 & dbs_latent_32_reg_segment_0);
  --mux write dbs 3, which is an e_mux
  descriptor_offset_bridge_m1_dbs_write_32 <= A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (internal_descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000000"))), descriptor_offset_bridge_m1_writedata(31 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (internal_descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000001"))), descriptor_offset_bridge_m1_writedata(63 DOWNTO 32), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (internal_descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000010"))), descriptor_offset_bridge_m1_writedata(95 DOWNTO 64), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (internal_descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000011"))), descriptor_offset_bridge_m1_writedata(127 DOWNTO 96), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (internal_descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000100"))), descriptor_offset_bridge_m1_writedata(159 DOWNTO 128), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (internal_descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000101"))), descriptor_offset_bridge_m1_writedata(191 DOWNTO 160), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (internal_descriptor_offset_bridge_m1_dbs_address(4 DOWNTO 2))) = std_logic_vector'("00000000000000000000000000000110"))), descriptor_offset_bridge_m1_writedata(223 DOWNTO 192), descriptor_offset_bridge_m1_writedata(255 DOWNTO 224))))))));
  --actual waitrequest port, which is an e_assign
  internal_descriptor_offset_bridge_m1_waitrequest <= NOT descriptor_offset_bridge_m1_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_descriptor_offset_bridge_m1_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_descriptor_offset_bridge_m1_latency_counter <= p1_descriptor_offset_bridge_m1_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_descriptor_offset_bridge_m1_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((descriptor_offset_bridge_m1_run AND ((descriptor_offset_bridge_m1_read AND descriptor_offset_bridge_m1_chipselect))))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_descriptor_offset_bridge_m1_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_descriptor_offset_bridge_m1_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_offset_bridge_m1_requests_descriptor_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --dbs count increment, which is an e_mux
  descriptor_offset_bridge_m1_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((descriptor_offset_bridge_m1_requests_descriptor_memory_s1)) = '1'), std_logic_vector'("00000000000000000000000000000100"), std_logic_vector'("00000000000000000000000000000000")), 5);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_descriptor_offset_bridge_m1_dbs_address(4) AND NOT((next_dbs_address(4)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_descriptor_offset_bridge_m1_dbs_address)) + (std_logic_vector'("0") & (descriptor_offset_bridge_m1_dbs_increment))), 5);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_descriptor_offset_bridge_m1_dbs_address <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_descriptor_offset_bridge_m1_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  descriptor_offset_bridge_m1_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (descriptor_offset_bridge_m1_dbs_rdv_counter)) + (std_logic_vector'("0") & (descriptor_offset_bridge_m1_dbs_rdv_counter_inc))), 5);
  --descriptor_offset_bridge_m1_rdv_inc_mux, which is an e_mux
  descriptor_offset_bridge_m1_dbs_rdv_counter_inc <= std_logic_vector'("00100");
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_offset_bridge_m1_dbs_rdv_counter <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        descriptor_offset_bridge_m1_dbs_rdv_counter <= descriptor_offset_bridge_m1_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= descriptor_offset_bridge_m1_dbs_rdv_counter(4) AND NOT descriptor_offset_bridge_m1_next_dbs_rdv_counter(4);
  --vhdl renameroo for output signals
  descriptor_offset_bridge_m1_address_to_slave <= internal_descriptor_offset_bridge_m1_address_to_slave;
  --vhdl renameroo for output signals
  descriptor_offset_bridge_m1_dbs_address <= internal_descriptor_offset_bridge_m1_dbs_address;
  --vhdl renameroo for output signals
  descriptor_offset_bridge_m1_latency_counter <= internal_descriptor_offset_bridge_m1_latency_counter;
  --vhdl renameroo for output signals
  descriptor_offset_bridge_m1_waitrequest <= internal_descriptor_offset_bridge_m1_waitrequest;
--synthesis translate_off
    --descriptor_offset_bridge_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        descriptor_offset_bridge_m1_address_last_time <= std_logic_vector'("000000000000000000000000000");
      elsif clk'event and clk = '1' then
        descriptor_offset_bridge_m1_address_last_time <= descriptor_offset_bridge_m1_address;
      end if;

    end process;

    --descriptor_offset_bridge/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_descriptor_offset_bridge_m1_waitrequest AND descriptor_offset_bridge_m1_chipselect;
      end if;

    end process;

    --descriptor_offset_bridge_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line18 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((descriptor_offset_bridge_m1_address /= descriptor_offset_bridge_m1_address_last_time))))) = '1' then 
          write(write_line18, now);
          write(write_line18, string'(": "));
          write(write_line18, string'("descriptor_offset_bridge_m1_address did not heed wait!!!"));
          write(output, write_line18.all);
          deallocate (write_line18);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --descriptor_offset_bridge_m1_chipselect check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        descriptor_offset_bridge_m1_chipselect_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        descriptor_offset_bridge_m1_chipselect_last_time <= descriptor_offset_bridge_m1_chipselect;
      end if;

    end process;

    --descriptor_offset_bridge_m1_chipselect matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line19 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(descriptor_offset_bridge_m1_chipselect) /= std_logic'(descriptor_offset_bridge_m1_chipselect_last_time)))))) = '1' then 
          write(write_line19, now);
          write(write_line19, string'(": "));
          write(write_line19, string'("descriptor_offset_bridge_m1_chipselect did not heed wait!!!"));
          write(output, write_line19.all);
          deallocate (write_line19);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --descriptor_offset_bridge_m1_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        descriptor_offset_bridge_m1_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        descriptor_offset_bridge_m1_burstcount_last_time <= descriptor_offset_bridge_m1_burstcount;
      end if;

    end process;

    --descriptor_offset_bridge_m1_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line20 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(descriptor_offset_bridge_m1_burstcount) /= std_logic'(descriptor_offset_bridge_m1_burstcount_last_time)))))) = '1' then 
          write(write_line20, now);
          write(write_line20, string'(": "));
          write(write_line20, string'("descriptor_offset_bridge_m1_burstcount did not heed wait!!!"));
          write(output, write_line20.all);
          deallocate (write_line20);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --descriptor_offset_bridge_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        descriptor_offset_bridge_m1_byteenable_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        descriptor_offset_bridge_m1_byteenable_last_time <= descriptor_offset_bridge_m1_byteenable;
      end if;

    end process;

    --descriptor_offset_bridge_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line21 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((descriptor_offset_bridge_m1_byteenable /= descriptor_offset_bridge_m1_byteenable_last_time))))) = '1' then 
          write(write_line21, now);
          write(write_line21, string'(": "));
          write(write_line21, string'("descriptor_offset_bridge_m1_byteenable did not heed wait!!!"));
          write(output, write_line21.all);
          deallocate (write_line21);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --descriptor_offset_bridge_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        descriptor_offset_bridge_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        descriptor_offset_bridge_m1_read_last_time <= descriptor_offset_bridge_m1_read;
      end if;

    end process;

    --descriptor_offset_bridge_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line22 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(descriptor_offset_bridge_m1_read) /= std_logic'(descriptor_offset_bridge_m1_read_last_time)))))) = '1' then 
          write(write_line22, now);
          write(write_line22, string'(": "));
          write(write_line22, string'("descriptor_offset_bridge_m1_read did not heed wait!!!"));
          write(output, write_line22.all);
          deallocate (write_line22);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --descriptor_offset_bridge_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        descriptor_offset_bridge_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        descriptor_offset_bridge_m1_write_last_time <= descriptor_offset_bridge_m1_write;
      end if;

    end process;

    --descriptor_offset_bridge_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line23 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(descriptor_offset_bridge_m1_write) /= std_logic'(descriptor_offset_bridge_m1_write_last_time)))))) = '1' then 
          write(write_line23, now);
          write(write_line23, string'(": "));
          write(write_line23, string'("descriptor_offset_bridge_m1_write did not heed wait!!!"));
          write(output, write_line23.all);
          deallocate (write_line23);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --descriptor_offset_bridge_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        descriptor_offset_bridge_m1_writedata_last_time <= std_logic_vector'("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        descriptor_offset_bridge_m1_writedata_last_time <= descriptor_offset_bridge_m1_writedata;
      end if;

    end process;

    --descriptor_offset_bridge_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line24 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((descriptor_offset_bridge_m1_writedata /= descriptor_offset_bridge_m1_writedata_last_time)))) AND ((descriptor_offset_bridge_m1_write AND descriptor_offset_bridge_m1_chipselect)))) = '1' then 
          write(write_line24, now);
          write(write_line24, string'(": "));
          write(write_line24, string'("descriptor_offset_bridge_m1_writedata did not heed wait!!!"));
          write(output, write_line24.all);
          deallocate (write_line24);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity descriptor_offset_bridge_bridge_arbitrator is 
end entity descriptor_offset_bridge_bridge_arbitrator;


architecture europa of descriptor_offset_bridge_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity fft_pipeline_0_avalon_slave_0_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal fft_pipeline_0_avalon_slave_0_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_fft_pipeline_0_avalon_slave_0 : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 : OUT STD_LOGIC;
                 signal d1_fft_pipeline_0_avalon_slave_0_end_xfer : OUT STD_LOGIC;
                 signal fft_pipeline_0_avalon_slave_0_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal fft_pipeline_0_avalon_slave_0_chipselect : OUT STD_LOGIC;
                 signal fft_pipeline_0_avalon_slave_0_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal fft_pipeline_0_avalon_slave_0_reset : OUT STD_LOGIC;
                 signal fft_pipeline_0_avalon_slave_0_write : OUT STD_LOGIC;
                 signal fft_pipeline_0_avalon_slave_0_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity fft_pipeline_0_avalon_slave_0_arbitrator;


architecture europa of fft_pipeline_0_avalon_slave_0_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_fft_pipeline_0_avalon_slave_0 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_fft_pipeline_0_avalon_slave_0 :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_allgrants :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_allow_new_arb_cycle :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_any_bursting_master_saved_grant :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_any_continuerequest :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_arb_counter_enable :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_arb_share_counter :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_arb_share_counter_next_value :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_arb_share_set_values :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_beginbursttransfer_internal :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_begins_xfer :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_end_xfer :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_firsttransfer :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_grant_vector :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_in_a_read_cycle :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_in_a_write_cycle :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_master_qreq_vector :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_non_bursting_master_requests :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_reg_firsttransfer :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_slavearbiterlockenable :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_slavearbiterlockenable2 :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_unreg_firsttransfer :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_waits_for_read :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 :  STD_LOGIC;
                signal shifted_address_to_fft_pipeline_0_avalon_slave_0_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_fft_pipeline_0_avalon_slave_0_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT fft_pipeline_0_avalon_slave_0_end_xfer;
    end if;

  end process;

  fft_pipeline_0_avalon_slave_0_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0);
  --assign fft_pipeline_0_avalon_slave_0_readdata_from_sa = fft_pipeline_0_avalon_slave_0_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  fft_pipeline_0_avalon_slave_0_readdata_from_sa <= fft_pipeline_0_avalon_slave_0_readdata;
  internal_cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("100000000000000000000000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --fft_pipeline_0_avalon_slave_0_arb_share_counter set values, which is an e_mux
  fft_pipeline_0_avalon_slave_0_arb_share_set_values <= std_logic'('1');
  --fft_pipeline_0_avalon_slave_0_non_bursting_master_requests mux, which is an e_mux
  fft_pipeline_0_avalon_slave_0_non_bursting_master_requests <= internal_cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0;
  --fft_pipeline_0_avalon_slave_0_any_bursting_master_saved_grant mux, which is an e_mux
  fft_pipeline_0_avalon_slave_0_any_bursting_master_saved_grant <= std_logic'('0');
  --fft_pipeline_0_avalon_slave_0_arb_share_counter_next_value assignment, which is an e_assign
  fft_pipeline_0_avalon_slave_0_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(fft_pipeline_0_avalon_slave_0_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(fft_pipeline_0_avalon_slave_0_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(fft_pipeline_0_avalon_slave_0_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(fft_pipeline_0_avalon_slave_0_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --fft_pipeline_0_avalon_slave_0_allgrants all slave grants, which is an e_mux
  fft_pipeline_0_avalon_slave_0_allgrants <= fft_pipeline_0_avalon_slave_0_grant_vector;
  --fft_pipeline_0_avalon_slave_0_end_xfer assignment, which is an e_assign
  fft_pipeline_0_avalon_slave_0_end_xfer <= NOT ((fft_pipeline_0_avalon_slave_0_waits_for_read OR fft_pipeline_0_avalon_slave_0_waits_for_write));
  --end_xfer_arb_share_counter_term_fft_pipeline_0_avalon_slave_0 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_fft_pipeline_0_avalon_slave_0 <= fft_pipeline_0_avalon_slave_0_end_xfer AND (((NOT fft_pipeline_0_avalon_slave_0_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --fft_pipeline_0_avalon_slave_0_arb_share_counter arbitration counter enable, which is an e_assign
  fft_pipeline_0_avalon_slave_0_arb_counter_enable <= ((end_xfer_arb_share_counter_term_fft_pipeline_0_avalon_slave_0 AND fft_pipeline_0_avalon_slave_0_allgrants)) OR ((end_xfer_arb_share_counter_term_fft_pipeline_0_avalon_slave_0 AND NOT fft_pipeline_0_avalon_slave_0_non_bursting_master_requests));
  --fft_pipeline_0_avalon_slave_0_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fft_pipeline_0_avalon_slave_0_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(fft_pipeline_0_avalon_slave_0_arb_counter_enable) = '1' then 
        fft_pipeline_0_avalon_slave_0_arb_share_counter <= fft_pipeline_0_avalon_slave_0_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --fft_pipeline_0_avalon_slave_0_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fft_pipeline_0_avalon_slave_0_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((fft_pipeline_0_avalon_slave_0_master_qreq_vector AND end_xfer_arb_share_counter_term_fft_pipeline_0_avalon_slave_0)) OR ((end_xfer_arb_share_counter_term_fft_pipeline_0_avalon_slave_0 AND NOT fft_pipeline_0_avalon_slave_0_non_bursting_master_requests)))) = '1' then 
        fft_pipeline_0_avalon_slave_0_slavearbiterlockenable <= fft_pipeline_0_avalon_slave_0_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master fft_pipeline_0/avalon_slave_0 arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= fft_pipeline_0_avalon_slave_0_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --fft_pipeline_0_avalon_slave_0_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  fft_pipeline_0_avalon_slave_0_slavearbiterlockenable2 <= fft_pipeline_0_avalon_slave_0_arb_share_counter_next_value;
  --cpuNios/data_master fft_pipeline_0/avalon_slave_0 arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= fft_pipeline_0_avalon_slave_0_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --fft_pipeline_0_avalon_slave_0_any_continuerequest at least one master continues requesting, which is an e_assign
  fft_pipeline_0_avalon_slave_0_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 <= internal_cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 AND NOT ((((cpuNios_data_master_read AND (NOT cpuNios_data_master_waitrequest))) OR (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write))));
  --fft_pipeline_0_avalon_slave_0_writedata mux, which is an e_mux
  fft_pipeline_0_avalon_slave_0_writedata <= cpuNios_data_master_writedata;
  --master is always granted when requested
  internal_cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 <= internal_cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0;
  --cpuNios/data_master saved-grant fft_pipeline_0/avalon_slave_0, which is an e_assign
  cpuNios_data_master_saved_grant_fft_pipeline_0_avalon_slave_0 <= internal_cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0;
  --allow new arb cycle for fft_pipeline_0/avalon_slave_0, which is an e_assign
  fft_pipeline_0_avalon_slave_0_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  fft_pipeline_0_avalon_slave_0_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  fft_pipeline_0_avalon_slave_0_master_qreq_vector <= std_logic'('1');
  --~fft_pipeline_0_avalon_slave_0_reset assignment, which is an e_assign
  fft_pipeline_0_avalon_slave_0_reset <= NOT reset_n;
  fft_pipeline_0_avalon_slave_0_chipselect <= internal_cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0;
  --fft_pipeline_0_avalon_slave_0_firsttransfer first transaction, which is an e_assign
  fft_pipeline_0_avalon_slave_0_firsttransfer <= A_WE_StdLogic((std_logic'(fft_pipeline_0_avalon_slave_0_begins_xfer) = '1'), fft_pipeline_0_avalon_slave_0_unreg_firsttransfer, fft_pipeline_0_avalon_slave_0_reg_firsttransfer);
  --fft_pipeline_0_avalon_slave_0_unreg_firsttransfer first transaction, which is an e_assign
  fft_pipeline_0_avalon_slave_0_unreg_firsttransfer <= NOT ((fft_pipeline_0_avalon_slave_0_slavearbiterlockenable AND fft_pipeline_0_avalon_slave_0_any_continuerequest));
  --fft_pipeline_0_avalon_slave_0_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fft_pipeline_0_avalon_slave_0_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(fft_pipeline_0_avalon_slave_0_begins_xfer) = '1' then 
        fft_pipeline_0_avalon_slave_0_reg_firsttransfer <= fft_pipeline_0_avalon_slave_0_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --fft_pipeline_0_avalon_slave_0_beginbursttransfer_internal begin burst transfer, which is an e_assign
  fft_pipeline_0_avalon_slave_0_beginbursttransfer_internal <= fft_pipeline_0_avalon_slave_0_begins_xfer;
  --fft_pipeline_0_avalon_slave_0_write assignment, which is an e_mux
  fft_pipeline_0_avalon_slave_0_write <= internal_cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 AND cpuNios_data_master_write;
  shifted_address_to_fft_pipeline_0_avalon_slave_0_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --fft_pipeline_0_avalon_slave_0_address mux, which is an e_mux
  fft_pipeline_0_avalon_slave_0_address <= A_EXT (A_SRL(shifted_address_to_fft_pipeline_0_avalon_slave_0_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")), 11);
  --d1_fft_pipeline_0_avalon_slave_0_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_fft_pipeline_0_avalon_slave_0_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_fft_pipeline_0_avalon_slave_0_end_xfer <= fft_pipeline_0_avalon_slave_0_end_xfer;
    end if;

  end process;

  --fft_pipeline_0_avalon_slave_0_waits_for_read in a cycle, which is an e_mux
  fft_pipeline_0_avalon_slave_0_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(fft_pipeline_0_avalon_slave_0_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --fft_pipeline_0_avalon_slave_0_in_a_read_cycle assignment, which is an e_assign
  fft_pipeline_0_avalon_slave_0_in_a_read_cycle <= internal_cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= fft_pipeline_0_avalon_slave_0_in_a_read_cycle;
  --fft_pipeline_0_avalon_slave_0_waits_for_write in a cycle, which is an e_mux
  fft_pipeline_0_avalon_slave_0_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(fft_pipeline_0_avalon_slave_0_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --fft_pipeline_0_avalon_slave_0_in_a_write_cycle assignment, which is an e_assign
  fft_pipeline_0_avalon_slave_0_in_a_write_cycle <= internal_cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= fft_pipeline_0_avalon_slave_0_in_a_write_cycle;
  wait_for_fft_pipeline_0_avalon_slave_0_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 <= internal_cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 <= internal_cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 <= internal_cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0;
--synthesis translate_off
    --fft_pipeline_0/avalon_slave_0 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity jtag_uart_avalon_jtag_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity jtag_uart_avalon_jtag_slave_arbitrator;


architecture europa of jtag_uart_avalon_jtag_slave_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allgrants :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_continuerequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_counter_enable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_counter :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_set_values :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_begins_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_grant_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_read_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_write_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_master_qreq_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_non_bursting_master_requests :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_unreg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_read :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_jtag_uart_avalon_jtag_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  jtag_uart_avalon_jtag_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave);
  --assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readdata_from_sa <= jtag_uart_avalon_jtag_slave_readdata;
  internal_cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("100000000000100100010000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_dataavailable_from_sa <= jtag_uart_avalon_jtag_slave_dataavailable;
  --assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readyfordata_from_sa <= jtag_uart_avalon_jtag_slave_readyfordata;
  --assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= jtag_uart_avalon_jtag_slave_waitrequest;
  --jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  jtag_uart_avalon_jtag_slave_arb_share_set_values <= std_logic'('1');
  --jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_non_bursting_master_requests <= internal_cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(jtag_uart_avalon_jtag_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_avalon_jtag_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(jtag_uart_avalon_jtag_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_avalon_jtag_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  jtag_uart_avalon_jtag_slave_allgrants <= jtag_uart_avalon_jtag_slave_grant_vector;
  --jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_end_xfer <= NOT ((jtag_uart_avalon_jtag_slave_waits_for_read OR jtag_uart_avalon_jtag_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave <= jtag_uart_avalon_jtag_slave_end_xfer AND (((NOT jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND jtag_uart_avalon_jtag_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests));
  --jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_arb_counter_enable) = '1' then 
        jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((jtag_uart_avalon_jtag_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests)))) = '1' then 
        jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
  --cpuNios/data_master jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  jtag_uart_avalon_jtag_slave_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave <= internal_cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave AND NOT ((((cpuNios_data_master_read AND (NOT cpuNios_data_master_waitrequest))) OR (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write))));
  --jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_writedata <= cpuNios_data_master_writedata;
  --master is always granted when requested
  internal_cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave <= internal_cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  --cpuNios/data_master saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  cpuNios_data_master_saved_grant_jtag_uart_avalon_jtag_slave <= internal_cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave;
  --allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  jtag_uart_avalon_jtag_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  jtag_uart_avalon_jtag_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  jtag_uart_avalon_jtag_slave_master_qreq_vector <= std_logic'('1');
  --jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_reset_n <= reset_n;
  jtag_uart_avalon_jtag_slave_chipselect <= internal_cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_firsttransfer <= A_WE_StdLogic((std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1'), jtag_uart_avalon_jtag_slave_unreg_firsttransfer, jtag_uart_avalon_jtag_slave_reg_firsttransfer);
  --jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_unreg_firsttransfer <= NOT ((jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND jtag_uart_avalon_jtag_slave_any_continuerequest));
  --jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1' then 
        jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  jtag_uart_avalon_jtag_slave_beginbursttransfer_internal <= jtag_uart_avalon_jtag_slave_begins_xfer;
  --~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_read_n <= NOT ((internal_cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave AND cpuNios_data_master_read));
  --~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_write_n <= NOT ((internal_cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave AND cpuNios_data_master_write));
  shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_jtag_uart_avalon_jtag_slave_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_read <= jtag_uart_avalon_jtag_slave_in_a_read_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_read_cycle <= internal_cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  --jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_write <= jtag_uart_avalon_jtag_slave_in_a_write_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_write_cycle <= internal_cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wait_for_jtag_uart_avalon_jtag_slave_counter <= std_logic'('0');
  --assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_irq_from_sa <= jtag_uart_avalon_jtag_slave_irq;
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave <= internal_cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave <= internal_cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave <= internal_cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
--synthesis translate_off
    --jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_24_to_8_bits_dfa_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_in_ready : IN STD_LOGIC;
                 signal lcd_pixel_converter_out_data : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal lcd_pixel_converter_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_pixel_converter_out_endofpacket : IN STD_LOGIC;
                 signal lcd_pixel_converter_out_startofpacket : IN STD_LOGIC;
                 signal lcd_pixel_converter_out_valid : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_24_to_8_bits_dfa_in_data : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal lcd_24_to_8_bits_dfa_in_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_24_to_8_bits_dfa_in_endofpacket : OUT STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_in_ready_from_sa : OUT STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_in_reset_n : OUT STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_in_startofpacket : OUT STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_in_valid : OUT STD_LOGIC
              );
end entity lcd_24_to_8_bits_dfa_in_arbitrator;


architecture europa of lcd_24_to_8_bits_dfa_in_arbitrator is

begin

  --mux lcd_24_to_8_bits_dfa_in_data, which is an e_mux
  lcd_24_to_8_bits_dfa_in_data <= lcd_pixel_converter_out_data;
  --mux lcd_24_to_8_bits_dfa_in_empty, which is an e_mux
  lcd_24_to_8_bits_dfa_in_empty <= lcd_pixel_converter_out_empty;
  --mux lcd_24_to_8_bits_dfa_in_endofpacket, which is an e_mux
  lcd_24_to_8_bits_dfa_in_endofpacket <= lcd_pixel_converter_out_endofpacket;
  --assign lcd_24_to_8_bits_dfa_in_ready_from_sa = lcd_24_to_8_bits_dfa_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_24_to_8_bits_dfa_in_ready_from_sa <= lcd_24_to_8_bits_dfa_in_ready;
  --mux lcd_24_to_8_bits_dfa_in_startofpacket, which is an e_mux
  lcd_24_to_8_bits_dfa_in_startofpacket <= lcd_pixel_converter_out_startofpacket;
  --mux lcd_24_to_8_bits_dfa_in_valid, which is an e_mux
  lcd_24_to_8_bits_dfa_in_valid <= lcd_pixel_converter_out_valid;
  --lcd_24_to_8_bits_dfa_in_reset_n assignment, which is an e_assign
  lcd_24_to_8_bits_dfa_in_reset_n <= reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_24_to_8_bits_dfa_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_out_data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal lcd_24_to_8_bits_dfa_out_empty : IN STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_out_endofpacket : IN STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_out_startofpacket : IN STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_out_valid : IN STD_LOGIC;
                 signal lcd_sync_generator_in_ready_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_24_to_8_bits_dfa_out_ready : OUT STD_LOGIC
              );
end entity lcd_24_to_8_bits_dfa_out_arbitrator;


architecture europa of lcd_24_to_8_bits_dfa_out_arbitrator is

begin

  --mux lcd_24_to_8_bits_dfa_out_ready, which is an e_mux
  lcd_24_to_8_bits_dfa_out_ready <= lcd_sync_generator_in_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_64_to_32_bits_dfa_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_in_ready : IN STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_ta_fifo_to_dfa_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_ta_fifo_to_dfa_out_endofpacket : IN STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_out_startofpacket : IN STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_out_valid : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_64_to_32_bits_dfa_in_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_64_to_32_bits_dfa_in_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_64_to_32_bits_dfa_in_endofpacket : OUT STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_in_ready_from_sa : OUT STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_in_reset_n : OUT STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_in_startofpacket : OUT STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_in_valid : OUT STD_LOGIC
              );
end entity lcd_64_to_32_bits_dfa_in_arbitrator;


architecture europa of lcd_64_to_32_bits_dfa_in_arbitrator is

begin

  --mux lcd_64_to_32_bits_dfa_in_data, which is an e_mux
  lcd_64_to_32_bits_dfa_in_data <= lcd_ta_fifo_to_dfa_out_data;
  --mux lcd_64_to_32_bits_dfa_in_empty, which is an e_mux
  lcd_64_to_32_bits_dfa_in_empty <= lcd_ta_fifo_to_dfa_out_empty;
  --mux lcd_64_to_32_bits_dfa_in_endofpacket, which is an e_mux
  lcd_64_to_32_bits_dfa_in_endofpacket <= lcd_ta_fifo_to_dfa_out_endofpacket;
  --assign lcd_64_to_32_bits_dfa_in_ready_from_sa = lcd_64_to_32_bits_dfa_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_64_to_32_bits_dfa_in_ready_from_sa <= lcd_64_to_32_bits_dfa_in_ready;
  --mux lcd_64_to_32_bits_dfa_in_startofpacket, which is an e_mux
  lcd_64_to_32_bits_dfa_in_startofpacket <= lcd_ta_fifo_to_dfa_out_startofpacket;
  --mux lcd_64_to_32_bits_dfa_in_valid, which is an e_mux
  lcd_64_to_32_bits_dfa_in_valid <= lcd_ta_fifo_to_dfa_out_valid;
  --lcd_64_to_32_bits_dfa_in_reset_n assignment, which is an e_assign
  lcd_64_to_32_bits_dfa_in_reset_n <= reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_64_to_32_bits_dfa_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_64_to_32_bits_dfa_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_64_to_32_bits_dfa_out_endofpacket : IN STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_out_startofpacket : IN STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_out_valid : IN STD_LOGIC;
                 signal lcd_pixel_converter_in_ready_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_64_to_32_bits_dfa_out_ready : OUT STD_LOGIC
              );
end entity lcd_64_to_32_bits_dfa_out_arbitrator;


architecture europa of lcd_64_to_32_bits_dfa_out_arbitrator is

begin

  --mux lcd_64_to_32_bits_dfa_out_ready, which is an e_mux
  lcd_64_to_32_bits_dfa_out_ready <= lcd_pixel_converter_in_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_i2c_en_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_i2c_en_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_granted_lcd_i2c_en_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_lcd_i2c_en_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_lcd_i2c_en_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_lcd_i2c_en_s1 : OUT STD_LOGIC;
                 signal d1_lcd_i2c_en_s1_end_xfer : OUT STD_LOGIC;
                 signal lcd_i2c_en_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_i2c_en_s1_chipselect : OUT STD_LOGIC;
                 signal lcd_i2c_en_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal lcd_i2c_en_s1_reset_n : OUT STD_LOGIC;
                 signal lcd_i2c_en_s1_write_n : OUT STD_LOGIC;
                 signal lcd_i2c_en_s1_writedata : OUT STD_LOGIC
              );
end entity lcd_i2c_en_s1_arbitrator;


architecture europa of lcd_i2c_en_s1_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_lcd_i2c_en_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_lcd_i2c_en_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_lcd_i2c_en_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_lcd_i2c_en_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_lcd_i2c_en_s1 :  STD_LOGIC;
                signal lcd_i2c_en_s1_allgrants :  STD_LOGIC;
                signal lcd_i2c_en_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal lcd_i2c_en_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal lcd_i2c_en_s1_any_continuerequest :  STD_LOGIC;
                signal lcd_i2c_en_s1_arb_counter_enable :  STD_LOGIC;
                signal lcd_i2c_en_s1_arb_share_counter :  STD_LOGIC;
                signal lcd_i2c_en_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal lcd_i2c_en_s1_arb_share_set_values :  STD_LOGIC;
                signal lcd_i2c_en_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal lcd_i2c_en_s1_begins_xfer :  STD_LOGIC;
                signal lcd_i2c_en_s1_end_xfer :  STD_LOGIC;
                signal lcd_i2c_en_s1_firsttransfer :  STD_LOGIC;
                signal lcd_i2c_en_s1_grant_vector :  STD_LOGIC;
                signal lcd_i2c_en_s1_in_a_read_cycle :  STD_LOGIC;
                signal lcd_i2c_en_s1_in_a_write_cycle :  STD_LOGIC;
                signal lcd_i2c_en_s1_master_qreq_vector :  STD_LOGIC;
                signal lcd_i2c_en_s1_non_bursting_master_requests :  STD_LOGIC;
                signal lcd_i2c_en_s1_reg_firsttransfer :  STD_LOGIC;
                signal lcd_i2c_en_s1_slavearbiterlockenable :  STD_LOGIC;
                signal lcd_i2c_en_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal lcd_i2c_en_s1_unreg_firsttransfer :  STD_LOGIC;
                signal lcd_i2c_en_s1_waits_for_read :  STD_LOGIC;
                signal lcd_i2c_en_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_lcd_i2c_en_s1_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_lcd_i2c_en_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT lcd_i2c_en_s1_end_xfer;
    end if;

  end process;

  lcd_i2c_en_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_lcd_i2c_en_s1);
  --assign lcd_i2c_en_s1_readdata_from_sa = lcd_i2c_en_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_i2c_en_s1_readdata_from_sa <= lcd_i2c_en_s1_readdata;
  internal_cpuNios_data_master_requests_lcd_i2c_en_s1 <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("100000000000100011110000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --lcd_i2c_en_s1_arb_share_counter set values, which is an e_mux
  lcd_i2c_en_s1_arb_share_set_values <= std_logic'('1');
  --lcd_i2c_en_s1_non_bursting_master_requests mux, which is an e_mux
  lcd_i2c_en_s1_non_bursting_master_requests <= internal_cpuNios_data_master_requests_lcd_i2c_en_s1;
  --lcd_i2c_en_s1_any_bursting_master_saved_grant mux, which is an e_mux
  lcd_i2c_en_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --lcd_i2c_en_s1_arb_share_counter_next_value assignment, which is an e_assign
  lcd_i2c_en_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(lcd_i2c_en_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_en_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(lcd_i2c_en_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_en_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --lcd_i2c_en_s1_allgrants all slave grants, which is an e_mux
  lcd_i2c_en_s1_allgrants <= lcd_i2c_en_s1_grant_vector;
  --lcd_i2c_en_s1_end_xfer assignment, which is an e_assign
  lcd_i2c_en_s1_end_xfer <= NOT ((lcd_i2c_en_s1_waits_for_read OR lcd_i2c_en_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_lcd_i2c_en_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_lcd_i2c_en_s1 <= lcd_i2c_en_s1_end_xfer AND (((NOT lcd_i2c_en_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --lcd_i2c_en_s1_arb_share_counter arbitration counter enable, which is an e_assign
  lcd_i2c_en_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_lcd_i2c_en_s1 AND lcd_i2c_en_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_lcd_i2c_en_s1 AND NOT lcd_i2c_en_s1_non_bursting_master_requests));
  --lcd_i2c_en_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_i2c_en_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_i2c_en_s1_arb_counter_enable) = '1' then 
        lcd_i2c_en_s1_arb_share_counter <= lcd_i2c_en_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --lcd_i2c_en_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_i2c_en_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((lcd_i2c_en_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_lcd_i2c_en_s1)) OR ((end_xfer_arb_share_counter_term_lcd_i2c_en_s1 AND NOT lcd_i2c_en_s1_non_bursting_master_requests)))) = '1' then 
        lcd_i2c_en_s1_slavearbiterlockenable <= lcd_i2c_en_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master lcd_i2c_en/s1 arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= lcd_i2c_en_s1_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --lcd_i2c_en_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  lcd_i2c_en_s1_slavearbiterlockenable2 <= lcd_i2c_en_s1_arb_share_counter_next_value;
  --cpuNios/data_master lcd_i2c_en/s1 arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= lcd_i2c_en_s1_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --lcd_i2c_en_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  lcd_i2c_en_s1_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_lcd_i2c_en_s1 <= internal_cpuNios_data_master_requests_lcd_i2c_en_s1 AND NOT (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write));
  --lcd_i2c_en_s1_writedata mux, which is an e_mux
  lcd_i2c_en_s1_writedata <= cpuNios_data_master_writedata(0);
  --master is always granted when requested
  internal_cpuNios_data_master_granted_lcd_i2c_en_s1 <= internal_cpuNios_data_master_qualified_request_lcd_i2c_en_s1;
  --cpuNios/data_master saved-grant lcd_i2c_en/s1, which is an e_assign
  cpuNios_data_master_saved_grant_lcd_i2c_en_s1 <= internal_cpuNios_data_master_requests_lcd_i2c_en_s1;
  --allow new arb cycle for lcd_i2c_en/s1, which is an e_assign
  lcd_i2c_en_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  lcd_i2c_en_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  lcd_i2c_en_s1_master_qreq_vector <= std_logic'('1');
  --lcd_i2c_en_s1_reset_n assignment, which is an e_assign
  lcd_i2c_en_s1_reset_n <= reset_n;
  lcd_i2c_en_s1_chipselect <= internal_cpuNios_data_master_granted_lcd_i2c_en_s1;
  --lcd_i2c_en_s1_firsttransfer first transaction, which is an e_assign
  lcd_i2c_en_s1_firsttransfer <= A_WE_StdLogic((std_logic'(lcd_i2c_en_s1_begins_xfer) = '1'), lcd_i2c_en_s1_unreg_firsttransfer, lcd_i2c_en_s1_reg_firsttransfer);
  --lcd_i2c_en_s1_unreg_firsttransfer first transaction, which is an e_assign
  lcd_i2c_en_s1_unreg_firsttransfer <= NOT ((lcd_i2c_en_s1_slavearbiterlockenable AND lcd_i2c_en_s1_any_continuerequest));
  --lcd_i2c_en_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_i2c_en_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_i2c_en_s1_begins_xfer) = '1' then 
        lcd_i2c_en_s1_reg_firsttransfer <= lcd_i2c_en_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --lcd_i2c_en_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  lcd_i2c_en_s1_beginbursttransfer_internal <= lcd_i2c_en_s1_begins_xfer;
  --~lcd_i2c_en_s1_write_n assignment, which is an e_mux
  lcd_i2c_en_s1_write_n <= NOT ((internal_cpuNios_data_master_granted_lcd_i2c_en_s1 AND cpuNios_data_master_write));
  shifted_address_to_lcd_i2c_en_s1_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --lcd_i2c_en_s1_address mux, which is an e_mux
  lcd_i2c_en_s1_address <= A_EXT (A_SRL(shifted_address_to_lcd_i2c_en_s1_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_lcd_i2c_en_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_lcd_i2c_en_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_lcd_i2c_en_s1_end_xfer <= lcd_i2c_en_s1_end_xfer;
    end if;

  end process;

  --lcd_i2c_en_s1_waits_for_read in a cycle, which is an e_mux
  lcd_i2c_en_s1_waits_for_read <= lcd_i2c_en_s1_in_a_read_cycle AND lcd_i2c_en_s1_begins_xfer;
  --lcd_i2c_en_s1_in_a_read_cycle assignment, which is an e_assign
  lcd_i2c_en_s1_in_a_read_cycle <= internal_cpuNios_data_master_granted_lcd_i2c_en_s1 AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= lcd_i2c_en_s1_in_a_read_cycle;
  --lcd_i2c_en_s1_waits_for_write in a cycle, which is an e_mux
  lcd_i2c_en_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_en_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --lcd_i2c_en_s1_in_a_write_cycle assignment, which is an e_assign
  lcd_i2c_en_s1_in_a_write_cycle <= internal_cpuNios_data_master_granted_lcd_i2c_en_s1 AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= lcd_i2c_en_s1_in_a_write_cycle;
  wait_for_lcd_i2c_en_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_lcd_i2c_en_s1 <= internal_cpuNios_data_master_granted_lcd_i2c_en_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_lcd_i2c_en_s1 <= internal_cpuNios_data_master_qualified_request_lcd_i2c_en_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_lcd_i2c_en_s1 <= internal_cpuNios_data_master_requests_lcd_i2c_en_s1;
--synthesis translate_off
    --lcd_i2c_en/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_i2c_scl_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_i2c_scl_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_granted_lcd_i2c_scl_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_lcd_i2c_scl_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_lcd_i2c_scl_s1 : OUT STD_LOGIC;
                 signal d1_lcd_i2c_scl_s1_end_xfer : OUT STD_LOGIC;
                 signal lcd_i2c_scl_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_i2c_scl_s1_chipselect : OUT STD_LOGIC;
                 signal lcd_i2c_scl_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal lcd_i2c_scl_s1_reset_n : OUT STD_LOGIC;
                 signal lcd_i2c_scl_s1_write_n : OUT STD_LOGIC;
                 signal lcd_i2c_scl_s1_writedata : OUT STD_LOGIC
              );
end entity lcd_i2c_scl_s1_arbitrator;


architecture europa of lcd_i2c_scl_s1_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_lcd_i2c_scl_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_lcd_i2c_scl_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_lcd_i2c_scl_s1 :  STD_LOGIC;
                signal lcd_i2c_scl_s1_allgrants :  STD_LOGIC;
                signal lcd_i2c_scl_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal lcd_i2c_scl_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal lcd_i2c_scl_s1_any_continuerequest :  STD_LOGIC;
                signal lcd_i2c_scl_s1_arb_counter_enable :  STD_LOGIC;
                signal lcd_i2c_scl_s1_arb_share_counter :  STD_LOGIC;
                signal lcd_i2c_scl_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal lcd_i2c_scl_s1_arb_share_set_values :  STD_LOGIC;
                signal lcd_i2c_scl_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal lcd_i2c_scl_s1_begins_xfer :  STD_LOGIC;
                signal lcd_i2c_scl_s1_end_xfer :  STD_LOGIC;
                signal lcd_i2c_scl_s1_firsttransfer :  STD_LOGIC;
                signal lcd_i2c_scl_s1_grant_vector :  STD_LOGIC;
                signal lcd_i2c_scl_s1_in_a_read_cycle :  STD_LOGIC;
                signal lcd_i2c_scl_s1_in_a_write_cycle :  STD_LOGIC;
                signal lcd_i2c_scl_s1_master_qreq_vector :  STD_LOGIC;
                signal lcd_i2c_scl_s1_non_bursting_master_requests :  STD_LOGIC;
                signal lcd_i2c_scl_s1_reg_firsttransfer :  STD_LOGIC;
                signal lcd_i2c_scl_s1_slavearbiterlockenable :  STD_LOGIC;
                signal lcd_i2c_scl_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal lcd_i2c_scl_s1_unreg_firsttransfer :  STD_LOGIC;
                signal lcd_i2c_scl_s1_waits_for_read :  STD_LOGIC;
                signal lcd_i2c_scl_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_lcd_i2c_scl_s1_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_lcd_i2c_scl_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT lcd_i2c_scl_s1_end_xfer;
    end if;

  end process;

  lcd_i2c_scl_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_lcd_i2c_scl_s1);
  --assign lcd_i2c_scl_s1_readdata_from_sa = lcd_i2c_scl_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_i2c_scl_s1_readdata_from_sa <= lcd_i2c_scl_s1_readdata;
  internal_cpuNios_data_master_requests_lcd_i2c_scl_s1 <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("100000000000100011100000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --lcd_i2c_scl_s1_arb_share_counter set values, which is an e_mux
  lcd_i2c_scl_s1_arb_share_set_values <= std_logic'('1');
  --lcd_i2c_scl_s1_non_bursting_master_requests mux, which is an e_mux
  lcd_i2c_scl_s1_non_bursting_master_requests <= internal_cpuNios_data_master_requests_lcd_i2c_scl_s1;
  --lcd_i2c_scl_s1_any_bursting_master_saved_grant mux, which is an e_mux
  lcd_i2c_scl_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --lcd_i2c_scl_s1_arb_share_counter_next_value assignment, which is an e_assign
  lcd_i2c_scl_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(lcd_i2c_scl_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_scl_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(lcd_i2c_scl_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_scl_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --lcd_i2c_scl_s1_allgrants all slave grants, which is an e_mux
  lcd_i2c_scl_s1_allgrants <= lcd_i2c_scl_s1_grant_vector;
  --lcd_i2c_scl_s1_end_xfer assignment, which is an e_assign
  lcd_i2c_scl_s1_end_xfer <= NOT ((lcd_i2c_scl_s1_waits_for_read OR lcd_i2c_scl_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 <= lcd_i2c_scl_s1_end_xfer AND (((NOT lcd_i2c_scl_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --lcd_i2c_scl_s1_arb_share_counter arbitration counter enable, which is an e_assign
  lcd_i2c_scl_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 AND lcd_i2c_scl_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 AND NOT lcd_i2c_scl_s1_non_bursting_master_requests));
  --lcd_i2c_scl_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_i2c_scl_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_i2c_scl_s1_arb_counter_enable) = '1' then 
        lcd_i2c_scl_s1_arb_share_counter <= lcd_i2c_scl_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --lcd_i2c_scl_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_i2c_scl_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((lcd_i2c_scl_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_lcd_i2c_scl_s1)) OR ((end_xfer_arb_share_counter_term_lcd_i2c_scl_s1 AND NOT lcd_i2c_scl_s1_non_bursting_master_requests)))) = '1' then 
        lcd_i2c_scl_s1_slavearbiterlockenable <= lcd_i2c_scl_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master lcd_i2c_scl/s1 arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= lcd_i2c_scl_s1_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --lcd_i2c_scl_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  lcd_i2c_scl_s1_slavearbiterlockenable2 <= lcd_i2c_scl_s1_arb_share_counter_next_value;
  --cpuNios/data_master lcd_i2c_scl/s1 arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= lcd_i2c_scl_s1_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --lcd_i2c_scl_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  lcd_i2c_scl_s1_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 <= internal_cpuNios_data_master_requests_lcd_i2c_scl_s1 AND NOT (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write));
  --lcd_i2c_scl_s1_writedata mux, which is an e_mux
  lcd_i2c_scl_s1_writedata <= cpuNios_data_master_writedata(0);
  --master is always granted when requested
  internal_cpuNios_data_master_granted_lcd_i2c_scl_s1 <= internal_cpuNios_data_master_qualified_request_lcd_i2c_scl_s1;
  --cpuNios/data_master saved-grant lcd_i2c_scl/s1, which is an e_assign
  cpuNios_data_master_saved_grant_lcd_i2c_scl_s1 <= internal_cpuNios_data_master_requests_lcd_i2c_scl_s1;
  --allow new arb cycle for lcd_i2c_scl/s1, which is an e_assign
  lcd_i2c_scl_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  lcd_i2c_scl_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  lcd_i2c_scl_s1_master_qreq_vector <= std_logic'('1');
  --lcd_i2c_scl_s1_reset_n assignment, which is an e_assign
  lcd_i2c_scl_s1_reset_n <= reset_n;
  lcd_i2c_scl_s1_chipselect <= internal_cpuNios_data_master_granted_lcd_i2c_scl_s1;
  --lcd_i2c_scl_s1_firsttransfer first transaction, which is an e_assign
  lcd_i2c_scl_s1_firsttransfer <= A_WE_StdLogic((std_logic'(lcd_i2c_scl_s1_begins_xfer) = '1'), lcd_i2c_scl_s1_unreg_firsttransfer, lcd_i2c_scl_s1_reg_firsttransfer);
  --lcd_i2c_scl_s1_unreg_firsttransfer first transaction, which is an e_assign
  lcd_i2c_scl_s1_unreg_firsttransfer <= NOT ((lcd_i2c_scl_s1_slavearbiterlockenable AND lcd_i2c_scl_s1_any_continuerequest));
  --lcd_i2c_scl_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_i2c_scl_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_i2c_scl_s1_begins_xfer) = '1' then 
        lcd_i2c_scl_s1_reg_firsttransfer <= lcd_i2c_scl_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --lcd_i2c_scl_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  lcd_i2c_scl_s1_beginbursttransfer_internal <= lcd_i2c_scl_s1_begins_xfer;
  --~lcd_i2c_scl_s1_write_n assignment, which is an e_mux
  lcd_i2c_scl_s1_write_n <= NOT ((internal_cpuNios_data_master_granted_lcd_i2c_scl_s1 AND cpuNios_data_master_write));
  shifted_address_to_lcd_i2c_scl_s1_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --lcd_i2c_scl_s1_address mux, which is an e_mux
  lcd_i2c_scl_s1_address <= A_EXT (A_SRL(shifted_address_to_lcd_i2c_scl_s1_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_lcd_i2c_scl_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_lcd_i2c_scl_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_lcd_i2c_scl_s1_end_xfer <= lcd_i2c_scl_s1_end_xfer;
    end if;

  end process;

  --lcd_i2c_scl_s1_waits_for_read in a cycle, which is an e_mux
  lcd_i2c_scl_s1_waits_for_read <= lcd_i2c_scl_s1_in_a_read_cycle AND lcd_i2c_scl_s1_begins_xfer;
  --lcd_i2c_scl_s1_in_a_read_cycle assignment, which is an e_assign
  lcd_i2c_scl_s1_in_a_read_cycle <= internal_cpuNios_data_master_granted_lcd_i2c_scl_s1 AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= lcd_i2c_scl_s1_in_a_read_cycle;
  --lcd_i2c_scl_s1_waits_for_write in a cycle, which is an e_mux
  lcd_i2c_scl_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_scl_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --lcd_i2c_scl_s1_in_a_write_cycle assignment, which is an e_assign
  lcd_i2c_scl_s1_in_a_write_cycle <= internal_cpuNios_data_master_granted_lcd_i2c_scl_s1 AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= lcd_i2c_scl_s1_in_a_write_cycle;
  wait_for_lcd_i2c_scl_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_lcd_i2c_scl_s1 <= internal_cpuNios_data_master_granted_lcd_i2c_scl_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 <= internal_cpuNios_data_master_qualified_request_lcd_i2c_scl_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_lcd_i2c_scl_s1 <= internal_cpuNios_data_master_requests_lcd_i2c_scl_s1;
--synthesis translate_off
    --lcd_i2c_scl/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_i2c_sdat_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_i2c_sdat_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_granted_lcd_i2c_sdat_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_lcd_i2c_sdat_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_lcd_i2c_sdat_s1 : OUT STD_LOGIC;
                 signal d1_lcd_i2c_sdat_s1_end_xfer : OUT STD_LOGIC;
                 signal lcd_i2c_sdat_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_i2c_sdat_s1_chipselect : OUT STD_LOGIC;
                 signal lcd_i2c_sdat_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal lcd_i2c_sdat_s1_reset_n : OUT STD_LOGIC;
                 signal lcd_i2c_sdat_s1_write_n : OUT STD_LOGIC;
                 signal lcd_i2c_sdat_s1_writedata : OUT STD_LOGIC
              );
end entity lcd_i2c_sdat_s1_arbitrator;


architecture europa of lcd_i2c_sdat_s1_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_lcd_i2c_sdat_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_lcd_i2c_sdat_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_lcd_i2c_sdat_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_lcd_i2c_sdat_s1 :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_allgrants :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_any_continuerequest :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_arb_counter_enable :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_arb_share_counter :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_arb_share_set_values :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_begins_xfer :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_end_xfer :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_firsttransfer :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_grant_vector :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_in_a_read_cycle :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_in_a_write_cycle :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_master_qreq_vector :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_non_bursting_master_requests :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_reg_firsttransfer :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_slavearbiterlockenable :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_unreg_firsttransfer :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_waits_for_read :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_lcd_i2c_sdat_s1_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_lcd_i2c_sdat_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT lcd_i2c_sdat_s1_end_xfer;
    end if;

  end process;

  lcd_i2c_sdat_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1);
  --assign lcd_i2c_sdat_s1_readdata_from_sa = lcd_i2c_sdat_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_i2c_sdat_s1_readdata_from_sa <= lcd_i2c_sdat_s1_readdata;
  internal_cpuNios_data_master_requests_lcd_i2c_sdat_s1 <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("100000000000100100000000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --lcd_i2c_sdat_s1_arb_share_counter set values, which is an e_mux
  lcd_i2c_sdat_s1_arb_share_set_values <= std_logic'('1');
  --lcd_i2c_sdat_s1_non_bursting_master_requests mux, which is an e_mux
  lcd_i2c_sdat_s1_non_bursting_master_requests <= internal_cpuNios_data_master_requests_lcd_i2c_sdat_s1;
  --lcd_i2c_sdat_s1_any_bursting_master_saved_grant mux, which is an e_mux
  lcd_i2c_sdat_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --lcd_i2c_sdat_s1_arb_share_counter_next_value assignment, which is an e_assign
  lcd_i2c_sdat_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(lcd_i2c_sdat_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_sdat_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(lcd_i2c_sdat_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_sdat_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --lcd_i2c_sdat_s1_allgrants all slave grants, which is an e_mux
  lcd_i2c_sdat_s1_allgrants <= lcd_i2c_sdat_s1_grant_vector;
  --lcd_i2c_sdat_s1_end_xfer assignment, which is an e_assign
  lcd_i2c_sdat_s1_end_xfer <= NOT ((lcd_i2c_sdat_s1_waits_for_read OR lcd_i2c_sdat_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_lcd_i2c_sdat_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_lcd_i2c_sdat_s1 <= lcd_i2c_sdat_s1_end_xfer AND (((NOT lcd_i2c_sdat_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --lcd_i2c_sdat_s1_arb_share_counter arbitration counter enable, which is an e_assign
  lcd_i2c_sdat_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_lcd_i2c_sdat_s1 AND lcd_i2c_sdat_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_lcd_i2c_sdat_s1 AND NOT lcd_i2c_sdat_s1_non_bursting_master_requests));
  --lcd_i2c_sdat_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_i2c_sdat_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_i2c_sdat_s1_arb_counter_enable) = '1' then 
        lcd_i2c_sdat_s1_arb_share_counter <= lcd_i2c_sdat_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --lcd_i2c_sdat_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_i2c_sdat_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((lcd_i2c_sdat_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_lcd_i2c_sdat_s1)) OR ((end_xfer_arb_share_counter_term_lcd_i2c_sdat_s1 AND NOT lcd_i2c_sdat_s1_non_bursting_master_requests)))) = '1' then 
        lcd_i2c_sdat_s1_slavearbiterlockenable <= lcd_i2c_sdat_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master lcd_i2c_sdat/s1 arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= lcd_i2c_sdat_s1_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --lcd_i2c_sdat_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  lcd_i2c_sdat_s1_slavearbiterlockenable2 <= lcd_i2c_sdat_s1_arb_share_counter_next_value;
  --cpuNios/data_master lcd_i2c_sdat/s1 arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= lcd_i2c_sdat_s1_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --lcd_i2c_sdat_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  lcd_i2c_sdat_s1_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 <= internal_cpuNios_data_master_requests_lcd_i2c_sdat_s1 AND NOT (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write));
  --lcd_i2c_sdat_s1_writedata mux, which is an e_mux
  lcd_i2c_sdat_s1_writedata <= cpuNios_data_master_writedata(0);
  --master is always granted when requested
  internal_cpuNios_data_master_granted_lcd_i2c_sdat_s1 <= internal_cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1;
  --cpuNios/data_master saved-grant lcd_i2c_sdat/s1, which is an e_assign
  cpuNios_data_master_saved_grant_lcd_i2c_sdat_s1 <= internal_cpuNios_data_master_requests_lcd_i2c_sdat_s1;
  --allow new arb cycle for lcd_i2c_sdat/s1, which is an e_assign
  lcd_i2c_sdat_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  lcd_i2c_sdat_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  lcd_i2c_sdat_s1_master_qreq_vector <= std_logic'('1');
  --lcd_i2c_sdat_s1_reset_n assignment, which is an e_assign
  lcd_i2c_sdat_s1_reset_n <= reset_n;
  lcd_i2c_sdat_s1_chipselect <= internal_cpuNios_data_master_granted_lcd_i2c_sdat_s1;
  --lcd_i2c_sdat_s1_firsttransfer first transaction, which is an e_assign
  lcd_i2c_sdat_s1_firsttransfer <= A_WE_StdLogic((std_logic'(lcd_i2c_sdat_s1_begins_xfer) = '1'), lcd_i2c_sdat_s1_unreg_firsttransfer, lcd_i2c_sdat_s1_reg_firsttransfer);
  --lcd_i2c_sdat_s1_unreg_firsttransfer first transaction, which is an e_assign
  lcd_i2c_sdat_s1_unreg_firsttransfer <= NOT ((lcd_i2c_sdat_s1_slavearbiterlockenable AND lcd_i2c_sdat_s1_any_continuerequest));
  --lcd_i2c_sdat_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_i2c_sdat_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_i2c_sdat_s1_begins_xfer) = '1' then 
        lcd_i2c_sdat_s1_reg_firsttransfer <= lcd_i2c_sdat_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --lcd_i2c_sdat_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  lcd_i2c_sdat_s1_beginbursttransfer_internal <= lcd_i2c_sdat_s1_begins_xfer;
  --~lcd_i2c_sdat_s1_write_n assignment, which is an e_mux
  lcd_i2c_sdat_s1_write_n <= NOT ((internal_cpuNios_data_master_granted_lcd_i2c_sdat_s1 AND cpuNios_data_master_write));
  shifted_address_to_lcd_i2c_sdat_s1_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --lcd_i2c_sdat_s1_address mux, which is an e_mux
  lcd_i2c_sdat_s1_address <= A_EXT (A_SRL(shifted_address_to_lcd_i2c_sdat_s1_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_lcd_i2c_sdat_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_lcd_i2c_sdat_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_lcd_i2c_sdat_s1_end_xfer <= lcd_i2c_sdat_s1_end_xfer;
    end if;

  end process;

  --lcd_i2c_sdat_s1_waits_for_read in a cycle, which is an e_mux
  lcd_i2c_sdat_s1_waits_for_read <= lcd_i2c_sdat_s1_in_a_read_cycle AND lcd_i2c_sdat_s1_begins_xfer;
  --lcd_i2c_sdat_s1_in_a_read_cycle assignment, which is an e_assign
  lcd_i2c_sdat_s1_in_a_read_cycle <= internal_cpuNios_data_master_granted_lcd_i2c_sdat_s1 AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= lcd_i2c_sdat_s1_in_a_read_cycle;
  --lcd_i2c_sdat_s1_waits_for_write in a cycle, which is an e_mux
  lcd_i2c_sdat_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_i2c_sdat_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --lcd_i2c_sdat_s1_in_a_write_cycle assignment, which is an e_assign
  lcd_i2c_sdat_s1_in_a_write_cycle <= internal_cpuNios_data_master_granted_lcd_i2c_sdat_s1 AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= lcd_i2c_sdat_s1_in_a_write_cycle;
  wait_for_lcd_i2c_sdat_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_lcd_i2c_sdat_s1 <= internal_cpuNios_data_master_granted_lcd_i2c_sdat_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 <= internal_cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_lcd_i2c_sdat_s1 <= internal_cpuNios_data_master_requests_lcd_i2c_sdat_s1;
--synthesis translate_off
    --lcd_i2c_sdat/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_pixel_converter_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_64_to_32_bits_dfa_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_64_to_32_bits_dfa_out_endofpacket : IN STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_out_startofpacket : IN STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_out_valid : IN STD_LOGIC;
                 signal lcd_pixel_converter_in_ready : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_pixel_converter_in_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_pixel_converter_in_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_pixel_converter_in_endofpacket : OUT STD_LOGIC;
                 signal lcd_pixel_converter_in_ready_from_sa : OUT STD_LOGIC;
                 signal lcd_pixel_converter_in_reset_n : OUT STD_LOGIC;
                 signal lcd_pixel_converter_in_startofpacket : OUT STD_LOGIC;
                 signal lcd_pixel_converter_in_valid : OUT STD_LOGIC
              );
end entity lcd_pixel_converter_in_arbitrator;


architecture europa of lcd_pixel_converter_in_arbitrator is

begin

  --mux lcd_pixel_converter_in_data, which is an e_mux
  lcd_pixel_converter_in_data <= lcd_64_to_32_bits_dfa_out_data;
  --mux lcd_pixel_converter_in_empty, which is an e_mux
  lcd_pixel_converter_in_empty <= lcd_64_to_32_bits_dfa_out_empty;
  --mux lcd_pixel_converter_in_endofpacket, which is an e_mux
  lcd_pixel_converter_in_endofpacket <= lcd_64_to_32_bits_dfa_out_endofpacket;
  --assign lcd_pixel_converter_in_ready_from_sa = lcd_pixel_converter_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_pixel_converter_in_ready_from_sa <= lcd_pixel_converter_in_ready;
  --mux lcd_pixel_converter_in_startofpacket, which is an e_mux
  lcd_pixel_converter_in_startofpacket <= lcd_64_to_32_bits_dfa_out_startofpacket;
  --mux lcd_pixel_converter_in_valid, which is an e_mux
  lcd_pixel_converter_in_valid <= lcd_64_to_32_bits_dfa_out_valid;
  --lcd_pixel_converter_in_reset_n assignment, which is an e_assign
  lcd_pixel_converter_in_reset_n <= reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_pixel_converter_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_in_ready_from_sa : IN STD_LOGIC;
                 signal lcd_pixel_converter_out_data : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal lcd_pixel_converter_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_pixel_converter_out_endofpacket : IN STD_LOGIC;
                 signal lcd_pixel_converter_out_startofpacket : IN STD_LOGIC;
                 signal lcd_pixel_converter_out_valid : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_pixel_converter_out_ready : OUT STD_LOGIC
              );
end entity lcd_pixel_converter_out_arbitrator;


architecture europa of lcd_pixel_converter_out_arbitrator is

begin

  --mux lcd_pixel_converter_out_ready, which is an e_mux
  lcd_pixel_converter_out_ready <= lcd_24_to_8_bits_dfa_in_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_pixel_fifo_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_pixel_fifo_in_ready : IN STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_ta_sgdma_to_fifo_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_ta_sgdma_to_fifo_out_endofpacket : IN STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_out_startofpacket : IN STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_out_valid : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_pixel_fifo_in_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_pixel_fifo_in_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_pixel_fifo_in_endofpacket : OUT STD_LOGIC;
                 signal lcd_pixel_fifo_in_ready_from_sa : OUT STD_LOGIC;
                 signal lcd_pixel_fifo_in_reset_n : OUT STD_LOGIC;
                 signal lcd_pixel_fifo_in_startofpacket : OUT STD_LOGIC;
                 signal lcd_pixel_fifo_in_valid : OUT STD_LOGIC
              );
end entity lcd_pixel_fifo_in_arbitrator;


architecture europa of lcd_pixel_fifo_in_arbitrator is

begin

  --mux lcd_pixel_fifo_in_data, which is an e_mux
  lcd_pixel_fifo_in_data <= lcd_ta_sgdma_to_fifo_out_data;
  --mux lcd_pixel_fifo_in_empty, which is an e_mux
  lcd_pixel_fifo_in_empty <= lcd_ta_sgdma_to_fifo_out_empty;
  --mux lcd_pixel_fifo_in_endofpacket, which is an e_mux
  lcd_pixel_fifo_in_endofpacket <= lcd_ta_sgdma_to_fifo_out_endofpacket;
  --assign lcd_pixel_fifo_in_ready_from_sa = lcd_pixel_fifo_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_pixel_fifo_in_ready_from_sa <= lcd_pixel_fifo_in_ready;
  --mux lcd_pixel_fifo_in_startofpacket, which is an e_mux
  lcd_pixel_fifo_in_startofpacket <= lcd_ta_sgdma_to_fifo_out_startofpacket;
  --mux lcd_pixel_fifo_in_valid, which is an e_mux
  lcd_pixel_fifo_in_valid <= lcd_ta_sgdma_to_fifo_out_valid;
  --lcd_pixel_fifo_in_reset_n assignment, which is an e_assign
  lcd_pixel_fifo_in_reset_n <= reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_pixel_fifo_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_pixel_fifo_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_pixel_fifo_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_pixel_fifo_out_endofpacket : IN STD_LOGIC;
                 signal lcd_pixel_fifo_out_startofpacket : IN STD_LOGIC;
                 signal lcd_pixel_fifo_out_valid : IN STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_in_ready_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_pixel_fifo_out_ready : OUT STD_LOGIC;
                 signal lcd_pixel_fifo_out_reset_n : OUT STD_LOGIC
              );
end entity lcd_pixel_fifo_out_arbitrator;


architecture europa of lcd_pixel_fifo_out_arbitrator is

begin

  --lcd_pixel_fifo_out_reset_n assignment, which is an e_assign
  lcd_pixel_fifo_out_reset_n <= reset_n;
  --mux lcd_pixel_fifo_out_ready, which is an e_mux
  lcd_pixel_fifo_out_ready <= lcd_ta_fifo_to_dfa_in_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_sgdma_csr_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_csr_irq : IN STD_LOGIC;
                 signal lcd_sgdma_csr_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr : OUT STD_LOGIC;
                 signal d1_lcd_sgdma_csr_end_xfer : OUT STD_LOGIC;
                 signal lcd_sgdma_csr_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal lcd_sgdma_csr_chipselect : OUT STD_LOGIC;
                 signal lcd_sgdma_csr_irq_from_sa : OUT STD_LOGIC;
                 signal lcd_sgdma_csr_read : OUT STD_LOGIC;
                 signal lcd_sgdma_csr_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_csr_reset_n : OUT STD_LOGIC;
                 signal lcd_sgdma_csr_write : OUT STD_LOGIC;
                 signal lcd_sgdma_csr_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity lcd_sgdma_csr_arbitrator;


architecture europa of lcd_sgdma_csr_arbitrator is
                signal cpu_ddr_clock_bridge_m1_arbiterlock :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_continuerequest :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_saved_grant_lcd_sgdma_csr :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_lcd_sgdma_csr :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr :  STD_LOGIC;
                signal lcd_sgdma_csr_allgrants :  STD_LOGIC;
                signal lcd_sgdma_csr_allow_new_arb_cycle :  STD_LOGIC;
                signal lcd_sgdma_csr_any_bursting_master_saved_grant :  STD_LOGIC;
                signal lcd_sgdma_csr_any_continuerequest :  STD_LOGIC;
                signal lcd_sgdma_csr_arb_counter_enable :  STD_LOGIC;
                signal lcd_sgdma_csr_arb_share_counter :  STD_LOGIC;
                signal lcd_sgdma_csr_arb_share_counter_next_value :  STD_LOGIC;
                signal lcd_sgdma_csr_arb_share_set_values :  STD_LOGIC;
                signal lcd_sgdma_csr_beginbursttransfer_internal :  STD_LOGIC;
                signal lcd_sgdma_csr_begins_xfer :  STD_LOGIC;
                signal lcd_sgdma_csr_end_xfer :  STD_LOGIC;
                signal lcd_sgdma_csr_firsttransfer :  STD_LOGIC;
                signal lcd_sgdma_csr_grant_vector :  STD_LOGIC;
                signal lcd_sgdma_csr_in_a_read_cycle :  STD_LOGIC;
                signal lcd_sgdma_csr_in_a_write_cycle :  STD_LOGIC;
                signal lcd_sgdma_csr_master_qreq_vector :  STD_LOGIC;
                signal lcd_sgdma_csr_non_bursting_master_requests :  STD_LOGIC;
                signal lcd_sgdma_csr_reg_firsttransfer :  STD_LOGIC;
                signal lcd_sgdma_csr_slavearbiterlockenable :  STD_LOGIC;
                signal lcd_sgdma_csr_slavearbiterlockenable2 :  STD_LOGIC;
                signal lcd_sgdma_csr_unreg_firsttransfer :  STD_LOGIC;
                signal lcd_sgdma_csr_waits_for_read :  STD_LOGIC;
                signal lcd_sgdma_csr_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_lcd_sgdma_csr_from_cpu_ddr_clock_bridge_m1 :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_lcd_sgdma_csr_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT lcd_sgdma_csr_end_xfer;
    end if;

  end process;

  lcd_sgdma_csr_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr);
  --assign lcd_sgdma_csr_readdata_from_sa = lcd_sgdma_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_sgdma_csr_readdata_from_sa <= lcd_sgdma_csr_readdata;
  internal_cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr <= to_std_logic(((Std_Logic_Vector'(cpu_ddr_clock_bridge_m1_address_to_slave(25 DOWNTO 6) & std_logic_vector'("000000")) = std_logic_vector'("10000000000000000000000000")))) AND ((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write));
  --lcd_sgdma_csr_arb_share_counter set values, which is an e_mux
  lcd_sgdma_csr_arb_share_set_values <= std_logic'('1');
  --lcd_sgdma_csr_non_bursting_master_requests mux, which is an e_mux
  lcd_sgdma_csr_non_bursting_master_requests <= internal_cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr;
  --lcd_sgdma_csr_any_bursting_master_saved_grant mux, which is an e_mux
  lcd_sgdma_csr_any_bursting_master_saved_grant <= std_logic'('0');
  --lcd_sgdma_csr_arb_share_counter_next_value assignment, which is an e_assign
  lcd_sgdma_csr_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(lcd_sgdma_csr_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_sgdma_csr_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(lcd_sgdma_csr_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_sgdma_csr_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --lcd_sgdma_csr_allgrants all slave grants, which is an e_mux
  lcd_sgdma_csr_allgrants <= lcd_sgdma_csr_grant_vector;
  --lcd_sgdma_csr_end_xfer assignment, which is an e_assign
  lcd_sgdma_csr_end_xfer <= NOT ((lcd_sgdma_csr_waits_for_read OR lcd_sgdma_csr_waits_for_write));
  --end_xfer_arb_share_counter_term_lcd_sgdma_csr arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_lcd_sgdma_csr <= lcd_sgdma_csr_end_xfer AND (((NOT lcd_sgdma_csr_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --lcd_sgdma_csr_arb_share_counter arbitration counter enable, which is an e_assign
  lcd_sgdma_csr_arb_counter_enable <= ((end_xfer_arb_share_counter_term_lcd_sgdma_csr AND lcd_sgdma_csr_allgrants)) OR ((end_xfer_arb_share_counter_term_lcd_sgdma_csr AND NOT lcd_sgdma_csr_non_bursting_master_requests));
  --lcd_sgdma_csr_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_sgdma_csr_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_sgdma_csr_arb_counter_enable) = '1' then 
        lcd_sgdma_csr_arb_share_counter <= lcd_sgdma_csr_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --lcd_sgdma_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_sgdma_csr_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((lcd_sgdma_csr_master_qreq_vector AND end_xfer_arb_share_counter_term_lcd_sgdma_csr)) OR ((end_xfer_arb_share_counter_term_lcd_sgdma_csr AND NOT lcd_sgdma_csr_non_bursting_master_requests)))) = '1' then 
        lcd_sgdma_csr_slavearbiterlockenable <= lcd_sgdma_csr_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_ddr_clock_bridge/m1 lcd_sgdma/csr arbiterlock, which is an e_assign
  cpu_ddr_clock_bridge_m1_arbiterlock <= lcd_sgdma_csr_slavearbiterlockenable AND cpu_ddr_clock_bridge_m1_continuerequest;
  --lcd_sgdma_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  lcd_sgdma_csr_slavearbiterlockenable2 <= lcd_sgdma_csr_arb_share_counter_next_value;
  --cpu_ddr_clock_bridge/m1 lcd_sgdma/csr arbiterlock2, which is an e_assign
  cpu_ddr_clock_bridge_m1_arbiterlock2 <= lcd_sgdma_csr_slavearbiterlockenable2 AND cpu_ddr_clock_bridge_m1_continuerequest;
  --lcd_sgdma_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  lcd_sgdma_csr_any_continuerequest <= std_logic'('1');
  --cpu_ddr_clock_bridge_m1_continuerequest continued request, which is an e_assign
  cpu_ddr_clock_bridge_m1_continuerequest <= std_logic'('1');
  internal_cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr <= internal_cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr AND NOT ((cpu_ddr_clock_bridge_m1_read AND ((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))) OR (cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register)))));
  --local readdatavalid cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr, which is an e_mux
  cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr <= (internal_cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr AND cpu_ddr_clock_bridge_m1_read) AND NOT lcd_sgdma_csr_waits_for_read;
  --lcd_sgdma_csr_writedata mux, which is an e_mux
  lcd_sgdma_csr_writedata <= cpu_ddr_clock_bridge_m1_writedata;
  --master is always granted when requested
  internal_cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr <= internal_cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr;
  --cpu_ddr_clock_bridge/m1 saved-grant lcd_sgdma/csr, which is an e_assign
  cpu_ddr_clock_bridge_m1_saved_grant_lcd_sgdma_csr <= internal_cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr;
  --allow new arb cycle for lcd_sgdma/csr, which is an e_assign
  lcd_sgdma_csr_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  lcd_sgdma_csr_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  lcd_sgdma_csr_master_qreq_vector <= std_logic'('1');
  --lcd_sgdma_csr_reset_n assignment, which is an e_assign
  lcd_sgdma_csr_reset_n <= reset_n;
  lcd_sgdma_csr_chipselect <= internal_cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr;
  --lcd_sgdma_csr_firsttransfer first transaction, which is an e_assign
  lcd_sgdma_csr_firsttransfer <= A_WE_StdLogic((std_logic'(lcd_sgdma_csr_begins_xfer) = '1'), lcd_sgdma_csr_unreg_firsttransfer, lcd_sgdma_csr_reg_firsttransfer);
  --lcd_sgdma_csr_unreg_firsttransfer first transaction, which is an e_assign
  lcd_sgdma_csr_unreg_firsttransfer <= NOT ((lcd_sgdma_csr_slavearbiterlockenable AND lcd_sgdma_csr_any_continuerequest));
  --lcd_sgdma_csr_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_sgdma_csr_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_sgdma_csr_begins_xfer) = '1' then 
        lcd_sgdma_csr_reg_firsttransfer <= lcd_sgdma_csr_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --lcd_sgdma_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  lcd_sgdma_csr_beginbursttransfer_internal <= lcd_sgdma_csr_begins_xfer;
  --lcd_sgdma_csr_read assignment, which is an e_mux
  lcd_sgdma_csr_read <= internal_cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr AND cpu_ddr_clock_bridge_m1_read;
  --lcd_sgdma_csr_write assignment, which is an e_mux
  lcd_sgdma_csr_write <= internal_cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr AND cpu_ddr_clock_bridge_m1_write;
  shifted_address_to_lcd_sgdma_csr_from_cpu_ddr_clock_bridge_m1 <= cpu_ddr_clock_bridge_m1_address_to_slave;
  --lcd_sgdma_csr_address mux, which is an e_mux
  lcd_sgdma_csr_address <= A_EXT (A_SRL(shifted_address_to_lcd_sgdma_csr_from_cpu_ddr_clock_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 4);
  --d1_lcd_sgdma_csr_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_lcd_sgdma_csr_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_lcd_sgdma_csr_end_xfer <= lcd_sgdma_csr_end_xfer;
    end if;

  end process;

  --lcd_sgdma_csr_waits_for_read in a cycle, which is an e_mux
  lcd_sgdma_csr_waits_for_read <= lcd_sgdma_csr_in_a_read_cycle AND lcd_sgdma_csr_begins_xfer;
  --lcd_sgdma_csr_in_a_read_cycle assignment, which is an e_assign
  lcd_sgdma_csr_in_a_read_cycle <= internal_cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr AND cpu_ddr_clock_bridge_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= lcd_sgdma_csr_in_a_read_cycle;
  --lcd_sgdma_csr_waits_for_write in a cycle, which is an e_mux
  lcd_sgdma_csr_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_sgdma_csr_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --lcd_sgdma_csr_in_a_write_cycle assignment, which is an e_assign
  lcd_sgdma_csr_in_a_write_cycle <= internal_cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr AND cpu_ddr_clock_bridge_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= lcd_sgdma_csr_in_a_write_cycle;
  wait_for_lcd_sgdma_csr_counter <= std_logic'('0');
  --assign lcd_sgdma_csr_irq_from_sa = lcd_sgdma_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_sgdma_csr_irq_from_sa <= lcd_sgdma_csr_irq;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr <= internal_cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr <= internal_cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr <= internal_cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr;
--synthesis translate_off
    --lcd_sgdma/csr enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_module;


architecture europa of selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity lcd_sgdma_descriptor_read_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_descriptor_read_granted_sdram_s1 : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_read : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_requests_sdram_s1 : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal lcd_sgdma_descriptor_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_descriptor_read_latency_counter : OUT STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_descriptor_read_readdatavalid : OUT STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_waitrequest : OUT STD_LOGIC
              );
end entity lcd_sgdma_descriptor_read_arbitrator;


architecture europa of lcd_sgdma_descriptor_read_arbitrator is
component selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_module;

                signal active_and_waiting_last_time :  STD_LOGIC;
                signal empty_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo :  STD_LOGIC;
                signal full_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo :  STD_LOGIC;
                signal internal_lcd_sgdma_descriptor_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_lcd_sgdma_descriptor_read_latency_counter :  STD_LOGIC;
                signal internal_lcd_sgdma_descriptor_read_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_descriptor_read_is_granted_some_slave :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_read_but_no_slave_selected :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_read_last_time :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_run :  STD_LOGIC;
                signal module_input15 :  STD_LOGIC;
                signal module_input16 :  STD_LOGIC;
                signal module_input17 :  STD_LOGIC;
                signal p1_lcd_sgdma_descriptor_read_latency_counter :  STD_LOGIC;
                signal pre_flush_lcd_sgdma_descriptor_read_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal read_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo :  STD_LOGIC;
                signal sdram_s1_readdata_from_sa_part_selected_by_negative_dbs :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_output :  STD_LOGIC;
                signal selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_output_sdram_s1 :  STD_LOGIC;
                signal write_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((lcd_sgdma_descriptor_read_qualified_request_sdram_s1 OR NOT lcd_sgdma_descriptor_read_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((lcd_sgdma_descriptor_read_granted_sdram_s1 OR NOT lcd_sgdma_descriptor_read_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT lcd_sgdma_descriptor_read_qualified_request_sdram_s1 OR NOT (lcd_sgdma_descriptor_read_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((lcd_sgdma_descriptor_read_read))))))))));
  --cascaded wait assignment, which is an e_assign
  lcd_sgdma_descriptor_read_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_lcd_sgdma_descriptor_read_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000000") & lcd_sgdma_descriptor_read_address(24 DOWNTO 0));
  --lcd_sgdma_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_sgdma_descriptor_read_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      lcd_sgdma_descriptor_read_read_but_no_slave_selected <= (lcd_sgdma_descriptor_read_read AND lcd_sgdma_descriptor_read_run) AND NOT lcd_sgdma_descriptor_read_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  lcd_sgdma_descriptor_read_is_granted_some_slave <= lcd_sgdma_descriptor_read_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_lcd_sgdma_descriptor_read_readdatavalid <= lcd_sgdma_descriptor_read_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  lcd_sgdma_descriptor_read_readdatavalid <= lcd_sgdma_descriptor_read_read_but_no_slave_selected OR pre_flush_lcd_sgdma_descriptor_read_readdatavalid;
  --Negative Dynamic Bus-sizing mux.
  --this mux selects the correct half of the 
  --wide data coming from the slave sdram/s1 
  sdram_s1_readdata_from_sa_part_selected_by_negative_dbs <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_output_sdram_s1))) = std_logic_vector'("00000000000000000000000000000000"))), sdram_s1_readdata_from_sa(31 DOWNTO 0), sdram_s1_readdata_from_sa(63 DOWNTO 32));
  --read_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo fifo read, which is an e_mux
  read_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo <= lcd_sgdma_descriptor_read_read_data_valid_sdram_s1;
  --write_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo fifo write, which is an e_mux
  write_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo <= (lcd_sgdma_descriptor_read_read AND lcd_sgdma_descriptor_read_run) AND lcd_sgdma_descriptor_read_requests_sdram_s1;
  selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_output_sdram_s1 <= selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_output;
  --selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo, which is an e_fifo_with_registered_outputs
  selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo : selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_module
    port map(
      data_out => selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo_output,
      empty => empty_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo,
      fifo_contains_ones_n => open,
      full => full_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo,
      clear_fifo => module_input15,
      clk => clk,
      data_in => module_input16,
      read => read_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo,
      reset_n => reset_n,
      sync_reset => module_input17,
      write => write_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo
    );

  module_input15 <= std_logic'('0');
  module_input16 <= internal_lcd_sgdma_descriptor_read_address_to_slave(2);
  module_input17 <= std_logic'('0');

  --lcd_sgdma/descriptor_read readdata mux, which is an e_mux
  lcd_sgdma_descriptor_read_readdata <= sdram_s1_readdata_from_sa_part_selected_by_negative_dbs;
  --actual waitrequest port, which is an e_assign
  internal_lcd_sgdma_descriptor_read_waitrequest <= NOT lcd_sgdma_descriptor_read_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_lcd_sgdma_descriptor_read_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_lcd_sgdma_descriptor_read_latency_counter <= p1_lcd_sgdma_descriptor_read_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_lcd_sgdma_descriptor_read_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((lcd_sgdma_descriptor_read_run AND lcd_sgdma_descriptor_read_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_read_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_lcd_sgdma_descriptor_read_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_read_address_to_slave <= internal_lcd_sgdma_descriptor_read_address_to_slave;
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_read_latency_counter <= internal_lcd_sgdma_descriptor_read_latency_counter;
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_read_waitrequest <= internal_lcd_sgdma_descriptor_read_waitrequest;
--synthesis translate_off
    --lcd_sgdma_descriptor_read_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        lcd_sgdma_descriptor_read_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        lcd_sgdma_descriptor_read_address_last_time <= lcd_sgdma_descriptor_read_address;
      end if;

    end process;

    --lcd_sgdma/descriptor_read waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_lcd_sgdma_descriptor_read_waitrequest AND (lcd_sgdma_descriptor_read_read);
      end if;

    end process;

    --lcd_sgdma_descriptor_read_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line25 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((lcd_sgdma_descriptor_read_address /= lcd_sgdma_descriptor_read_address_last_time))))) = '1' then 
          write(write_line25, now);
          write(write_line25, string'(": "));
          write(write_line25, string'("lcd_sgdma_descriptor_read_address did not heed wait!!!"));
          write(output, write_line25.all);
          deallocate (write_line25);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --lcd_sgdma_descriptor_read_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        lcd_sgdma_descriptor_read_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        lcd_sgdma_descriptor_read_read_last_time <= lcd_sgdma_descriptor_read_read;
      end if;

    end process;

    --lcd_sgdma_descriptor_read_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line26 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(lcd_sgdma_descriptor_read_read) /= std_logic'(lcd_sgdma_descriptor_read_read_last_time)))))) = '1' then 
          write(write_line26, now);
          write(write_line26, string'(": "));
          write(write_line26, string'("lcd_sgdma_descriptor_read_read did not heed wait!!!"));
          write(output, write_line26.all);
          deallocate (write_line26);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo read when empty, which is an e_process
    process (clk)
    VARIABLE write_line27 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((empty_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo AND read_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo)) = '1' then 
          write(write_line27, now);
          write(write_line27, string'(": "));
          write(write_line27, string'("lcd_sgdma/descriptor_read negative rdv fifo selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo: read AND empty."));
          write(output, write_line27.all & CR);
          deallocate (write_line27);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo write when full, which is an e_process
    process (clk)
    VARIABLE write_line28 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((full_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo AND write_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo) AND NOT read_selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo)) = '1' then 
          write(write_line28, now);
          write(write_line28, string'(": "));
          write(write_line28, string'("lcd_sgdma/descriptor_read negative rdv fifo selecto_nrdv_lcd_sgdma_descriptor_read_1_sdram_s1_fifo: write AND full."));
          write(output, write_line28.all & CR);
          deallocate (write_line28);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity lcd_sgdma_descriptor_write_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_descriptor_write_granted_sdram_s1 : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_write_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_write_requests_sdram_s1 : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_write_write : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal lcd_sgdma_descriptor_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_descriptor_write_waitrequest : OUT STD_LOGIC
              );
end entity lcd_sgdma_descriptor_write_arbitrator;


architecture europa of lcd_sgdma_descriptor_write_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_lcd_sgdma_descriptor_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_lcd_sgdma_descriptor_write_waitrequest :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_descriptor_write_run :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_write_last_time :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((lcd_sgdma_descriptor_write_qualified_request_sdram_s1 OR NOT lcd_sgdma_descriptor_write_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((lcd_sgdma_descriptor_write_granted_sdram_s1 OR NOT lcd_sgdma_descriptor_write_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT lcd_sgdma_descriptor_write_qualified_request_sdram_s1 OR NOT (lcd_sgdma_descriptor_write_write))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((lcd_sgdma_descriptor_write_write))))))))));
  --cascaded wait assignment, which is an e_assign
  lcd_sgdma_descriptor_write_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_lcd_sgdma_descriptor_write_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000000") & lcd_sgdma_descriptor_write_address(24 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_lcd_sgdma_descriptor_write_waitrequest <= NOT lcd_sgdma_descriptor_write_run;
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_write_address_to_slave <= internal_lcd_sgdma_descriptor_write_address_to_slave;
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_write_waitrequest <= internal_lcd_sgdma_descriptor_write_waitrequest;
--synthesis translate_off
    --lcd_sgdma_descriptor_write_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        lcd_sgdma_descriptor_write_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        lcd_sgdma_descriptor_write_address_last_time <= lcd_sgdma_descriptor_write_address;
      end if;

    end process;

    --lcd_sgdma/descriptor_write waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_lcd_sgdma_descriptor_write_waitrequest AND (lcd_sgdma_descriptor_write_write);
      end if;

    end process;

    --lcd_sgdma_descriptor_write_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line29 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((lcd_sgdma_descriptor_write_address /= lcd_sgdma_descriptor_write_address_last_time))))) = '1' then 
          write(write_line29, now);
          write(write_line29, string'(": "));
          write(write_line29, string'("lcd_sgdma_descriptor_write_address did not heed wait!!!"));
          write(output, write_line29.all);
          deallocate (write_line29);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --lcd_sgdma_descriptor_write_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        lcd_sgdma_descriptor_write_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        lcd_sgdma_descriptor_write_write_last_time <= lcd_sgdma_descriptor_write_write;
      end if;

    end process;

    --lcd_sgdma_descriptor_write_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line30 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(lcd_sgdma_descriptor_write_write) /= std_logic'(lcd_sgdma_descriptor_write_write_last_time)))))) = '1' then 
          write(write_line30, now);
          write(write_line30, string'(": "));
          write(write_line30, string'("lcd_sgdma_descriptor_write_write did not heed wait!!!"));
          write(output, write_line30.all);
          deallocate (write_line30);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --lcd_sgdma_descriptor_write_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        lcd_sgdma_descriptor_write_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        lcd_sgdma_descriptor_write_writedata_last_time <= lcd_sgdma_descriptor_write_writedata;
      end if;

    end process;

    --lcd_sgdma_descriptor_write_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line31 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((lcd_sgdma_descriptor_write_writedata /= lcd_sgdma_descriptor_write_writedata_last_time)))) AND lcd_sgdma_descriptor_write_write)) = '1' then 
          write(write_line31, now);
          write(write_line31, string'(": "));
          write(write_line31, string'("lcd_sgdma_descriptor_write_writedata did not heed wait!!!"));
          write(output, write_line31.all);
          deallocate (write_line31);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity lcd_sgdma_m_read_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal lcd_sgdma_m_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_m_read_granted_sdram_s1 : IN STD_LOGIC;
                 signal lcd_sgdma_m_read_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal lcd_sgdma_m_read_read : IN STD_LOGIC;
                 signal lcd_sgdma_m_read_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal lcd_sgdma_m_read_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal lcd_sgdma_m_read_requests_sdram_s1 : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal lcd_sgdma_m_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_m_read_latency_counter : OUT STD_LOGIC;
                 signal lcd_sgdma_m_read_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_sgdma_m_read_readdatavalid : OUT STD_LOGIC;
                 signal lcd_sgdma_m_read_waitrequest : OUT STD_LOGIC
              );
end entity lcd_sgdma_m_read_arbitrator;


architecture europa of lcd_sgdma_m_read_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_lcd_sgdma_m_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_lcd_sgdma_m_read_latency_counter :  STD_LOGIC;
                signal internal_lcd_sgdma_m_read_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal lcd_sgdma_m_read_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_m_read_is_granted_some_slave :  STD_LOGIC;
                signal lcd_sgdma_m_read_read_but_no_slave_selected :  STD_LOGIC;
                signal lcd_sgdma_m_read_read_last_time :  STD_LOGIC;
                signal lcd_sgdma_m_read_run :  STD_LOGIC;
                signal p1_lcd_sgdma_m_read_latency_counter :  STD_LOGIC;
                signal pre_flush_lcd_sgdma_m_read_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((lcd_sgdma_m_read_qualified_request_sdram_s1 OR NOT lcd_sgdma_m_read_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((lcd_sgdma_m_read_granted_sdram_s1 OR NOT lcd_sgdma_m_read_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT lcd_sgdma_m_read_qualified_request_sdram_s1 OR NOT (lcd_sgdma_m_read_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((lcd_sgdma_m_read_read))))))))));
  --cascaded wait assignment, which is an e_assign
  lcd_sgdma_m_read_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_lcd_sgdma_m_read_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000000") & lcd_sgdma_m_read_address(24 DOWNTO 0));
  --lcd_sgdma_m_read_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_sgdma_m_read_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      lcd_sgdma_m_read_read_but_no_slave_selected <= (lcd_sgdma_m_read_read AND lcd_sgdma_m_read_run) AND NOT lcd_sgdma_m_read_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  lcd_sgdma_m_read_is_granted_some_slave <= lcd_sgdma_m_read_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_lcd_sgdma_m_read_readdatavalid <= lcd_sgdma_m_read_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  lcd_sgdma_m_read_readdatavalid <= lcd_sgdma_m_read_read_but_no_slave_selected OR pre_flush_lcd_sgdma_m_read_readdatavalid;
  --lcd_sgdma/m_read readdata mux, which is an e_mux
  lcd_sgdma_m_read_readdata <= sdram_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_lcd_sgdma_m_read_waitrequest <= NOT lcd_sgdma_m_read_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_lcd_sgdma_m_read_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_lcd_sgdma_m_read_latency_counter <= p1_lcd_sgdma_m_read_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_lcd_sgdma_m_read_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((lcd_sgdma_m_read_run AND lcd_sgdma_m_read_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_m_read_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_lcd_sgdma_m_read_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --vhdl renameroo for output signals
  lcd_sgdma_m_read_address_to_slave <= internal_lcd_sgdma_m_read_address_to_slave;
  --vhdl renameroo for output signals
  lcd_sgdma_m_read_latency_counter <= internal_lcd_sgdma_m_read_latency_counter;
  --vhdl renameroo for output signals
  lcd_sgdma_m_read_waitrequest <= internal_lcd_sgdma_m_read_waitrequest;
--synthesis translate_off
    --lcd_sgdma_m_read_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        lcd_sgdma_m_read_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        lcd_sgdma_m_read_address_last_time <= lcd_sgdma_m_read_address;
      end if;

    end process;

    --lcd_sgdma/m_read waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_lcd_sgdma_m_read_waitrequest AND (lcd_sgdma_m_read_read);
      end if;

    end process;

    --lcd_sgdma_m_read_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line32 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((lcd_sgdma_m_read_address /= lcd_sgdma_m_read_address_last_time))))) = '1' then 
          write(write_line32, now);
          write(write_line32, string'(": "));
          write(write_line32, string'("lcd_sgdma_m_read_address did not heed wait!!!"));
          write(output, write_line32.all);
          deallocate (write_line32);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --lcd_sgdma_m_read_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        lcd_sgdma_m_read_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        lcd_sgdma_m_read_read_last_time <= lcd_sgdma_m_read_read;
      end if;

    end process;

    --lcd_sgdma_m_read_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line33 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(lcd_sgdma_m_read_read) /= std_logic'(lcd_sgdma_m_read_read_last_time)))))) = '1' then 
          write(write_line33, now);
          write(write_line33, string'(": "));
          write(write_line33, string'("lcd_sgdma_m_read_read did not heed wait!!!"));
          write(output, write_line33.all);
          deallocate (write_line33);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_sgdma_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_sgdma_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_sgdma_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_sgdma_out_endofpacket : IN STD_LOGIC;
                 signal lcd_sgdma_out_startofpacket : IN STD_LOGIC;
                 signal lcd_sgdma_out_valid : IN STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_in_ready_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_sgdma_out_ready : OUT STD_LOGIC
              );
end entity lcd_sgdma_out_arbitrator;


architecture europa of lcd_sgdma_out_arbitrator is

begin

  --mux lcd_sgdma_out_ready, which is an e_mux
  lcd_sgdma_out_ready <= lcd_ta_sgdma_to_fifo_in_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_sync_generator_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_out_data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal lcd_24_to_8_bits_dfa_out_empty : IN STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_out_endofpacket : IN STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_out_startofpacket : IN STD_LOGIC;
                 signal lcd_24_to_8_bits_dfa_out_valid : IN STD_LOGIC;
                 signal lcd_sync_generator_in_ready : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_sync_generator_in_data : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal lcd_sync_generator_in_empty : OUT STD_LOGIC;
                 signal lcd_sync_generator_in_endofpacket : OUT STD_LOGIC;
                 signal lcd_sync_generator_in_ready_from_sa : OUT STD_LOGIC;
                 signal lcd_sync_generator_in_reset_n : OUT STD_LOGIC;
                 signal lcd_sync_generator_in_startofpacket : OUT STD_LOGIC;
                 signal lcd_sync_generator_in_valid : OUT STD_LOGIC
              );
end entity lcd_sync_generator_in_arbitrator;


architecture europa of lcd_sync_generator_in_arbitrator is

begin

  --mux lcd_sync_generator_in_data, which is an e_mux
  lcd_sync_generator_in_data <= lcd_24_to_8_bits_dfa_out_data;
  --mux lcd_sync_generator_in_empty, which is an e_mux
  lcd_sync_generator_in_empty <= lcd_24_to_8_bits_dfa_out_empty;
  --mux lcd_sync_generator_in_endofpacket, which is an e_mux
  lcd_sync_generator_in_endofpacket <= lcd_24_to_8_bits_dfa_out_endofpacket;
  --assign lcd_sync_generator_in_ready_from_sa = lcd_sync_generator_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_sync_generator_in_ready_from_sa <= lcd_sync_generator_in_ready;
  --mux lcd_sync_generator_in_startofpacket, which is an e_mux
  lcd_sync_generator_in_startofpacket <= lcd_24_to_8_bits_dfa_out_startofpacket;
  --mux lcd_sync_generator_in_valid, which is an e_mux
  lcd_sync_generator_in_valid <= lcd_24_to_8_bits_dfa_out_valid;
  --lcd_sync_generator_in_reset_n assignment, which is an e_assign
  lcd_sync_generator_in_reset_n <= reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_ta_fifo_to_dfa_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_pixel_fifo_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_pixel_fifo_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_pixel_fifo_out_endofpacket : IN STD_LOGIC;
                 signal lcd_pixel_fifo_out_startofpacket : IN STD_LOGIC;
                 signal lcd_pixel_fifo_out_valid : IN STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_in_ready : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_ta_fifo_to_dfa_in_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_ta_fifo_to_dfa_in_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_ta_fifo_to_dfa_in_endofpacket : OUT STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_in_ready_from_sa : OUT STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_in_reset_n : OUT STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_in_startofpacket : OUT STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_in_valid : OUT STD_LOGIC
              );
end entity lcd_ta_fifo_to_dfa_in_arbitrator;


architecture europa of lcd_ta_fifo_to_dfa_in_arbitrator is

begin

  --mux lcd_ta_fifo_to_dfa_in_data, which is an e_mux
  lcd_ta_fifo_to_dfa_in_data <= lcd_pixel_fifo_out_data;
  --mux lcd_ta_fifo_to_dfa_in_empty, which is an e_mux
  lcd_ta_fifo_to_dfa_in_empty <= lcd_pixel_fifo_out_empty;
  --mux lcd_ta_fifo_to_dfa_in_endofpacket, which is an e_mux
  lcd_ta_fifo_to_dfa_in_endofpacket <= lcd_pixel_fifo_out_endofpacket;
  --assign lcd_ta_fifo_to_dfa_in_ready_from_sa = lcd_ta_fifo_to_dfa_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_ta_fifo_to_dfa_in_ready_from_sa <= lcd_ta_fifo_to_dfa_in_ready;
  --mux lcd_ta_fifo_to_dfa_in_startofpacket, which is an e_mux
  lcd_ta_fifo_to_dfa_in_startofpacket <= lcd_pixel_fifo_out_startofpacket;
  --mux lcd_ta_fifo_to_dfa_in_valid, which is an e_mux
  lcd_ta_fifo_to_dfa_in_valid <= lcd_pixel_fifo_out_valid;
  --lcd_ta_fifo_to_dfa_in_reset_n assignment, which is an e_assign
  lcd_ta_fifo_to_dfa_in_reset_n <= reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_ta_fifo_to_dfa_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_64_to_32_bits_dfa_in_ready_from_sa : IN STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_ta_fifo_to_dfa_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_ta_fifo_to_dfa_out_endofpacket : IN STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_out_startofpacket : IN STD_LOGIC;
                 signal lcd_ta_fifo_to_dfa_out_valid : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_ta_fifo_to_dfa_out_ready : OUT STD_LOGIC
              );
end entity lcd_ta_fifo_to_dfa_out_arbitrator;


architecture europa of lcd_ta_fifo_to_dfa_out_arbitrator is

begin

  --mux lcd_ta_fifo_to_dfa_out_ready, which is an e_mux
  lcd_ta_fifo_to_dfa_out_ready <= lcd_64_to_32_bits_dfa_in_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_ta_sgdma_to_fifo_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_sgdma_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_sgdma_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_sgdma_out_endofpacket : IN STD_LOGIC;
                 signal lcd_sgdma_out_startofpacket : IN STD_LOGIC;
                 signal lcd_sgdma_out_valid : IN STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_in_ready : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_ta_sgdma_to_fifo_in_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_ta_sgdma_to_fifo_in_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_ta_sgdma_to_fifo_in_endofpacket : OUT STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_in_ready_from_sa : OUT STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_in_reset_n : OUT STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_in_startofpacket : OUT STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_in_valid : OUT STD_LOGIC
              );
end entity lcd_ta_sgdma_to_fifo_in_arbitrator;


architecture europa of lcd_ta_sgdma_to_fifo_in_arbitrator is

begin

  --mux lcd_ta_sgdma_to_fifo_in_data, which is an e_mux
  lcd_ta_sgdma_to_fifo_in_data <= lcd_sgdma_out_data;
  --mux lcd_ta_sgdma_to_fifo_in_empty, which is an e_mux
  lcd_ta_sgdma_to_fifo_in_empty <= lcd_sgdma_out_empty;
  --mux lcd_ta_sgdma_to_fifo_in_endofpacket, which is an e_mux
  lcd_ta_sgdma_to_fifo_in_endofpacket <= lcd_sgdma_out_endofpacket;
  --assign lcd_ta_sgdma_to_fifo_in_ready_from_sa = lcd_ta_sgdma_to_fifo_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_ta_sgdma_to_fifo_in_ready_from_sa <= lcd_ta_sgdma_to_fifo_in_ready;
  --mux lcd_ta_sgdma_to_fifo_in_startofpacket, which is an e_mux
  lcd_ta_sgdma_to_fifo_in_startofpacket <= lcd_sgdma_out_startofpacket;
  --mux lcd_ta_sgdma_to_fifo_in_valid, which is an e_mux
  lcd_ta_sgdma_to_fifo_in_valid <= lcd_sgdma_out_valid;
  --lcd_ta_sgdma_to_fifo_in_reset_n assignment, which is an e_assign
  lcd_ta_sgdma_to_fifo_in_reset_n <= reset_n;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lcd_ta_sgdma_to_fifo_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_pixel_fifo_in_ready_from_sa : IN STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal lcd_ta_sgdma_to_fifo_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal lcd_ta_sgdma_to_fifo_out_endofpacket : IN STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_out_startofpacket : IN STD_LOGIC;
                 signal lcd_ta_sgdma_to_fifo_out_valid : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal lcd_ta_sgdma_to_fifo_out_ready : OUT STD_LOGIC
              );
end entity lcd_ta_sgdma_to_fifo_out_arbitrator;


architecture europa of lcd_ta_sgdma_to_fifo_out_arbitrator is

begin

  --mux lcd_ta_sgdma_to_fifo_out_ready, which is an e_mux
  lcd_ta_sgdma_to_fifo_out_ready <= lcd_pixel_fifo_in_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity performance_counter_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal performance_counter_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_granted_performance_counter_control_slave : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_performance_counter_control_slave : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_performance_counter_control_slave : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_performance_counter_control_slave : OUT STD_LOGIC;
                 signal d1_performance_counter_control_slave_end_xfer : OUT STD_LOGIC;
                 signal performance_counter_control_slave_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal performance_counter_control_slave_begintransfer : OUT STD_LOGIC;
                 signal performance_counter_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal performance_counter_control_slave_reset_n : OUT STD_LOGIC;
                 signal performance_counter_control_slave_write : OUT STD_LOGIC;
                 signal performance_counter_control_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave : OUT STD_LOGIC
              );
end entity performance_counter_control_slave_arbitrator;


architecture europa of performance_counter_control_slave_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register_in :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_performance_counter_control_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_performance_counter_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_performance_counter_control_slave :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_performance_counter_control_slave :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_performance_counter_control_slave :  STD_LOGIC;
                signal p1_cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register :  STD_LOGIC;
                signal performance_counter_control_slave_allgrants :  STD_LOGIC;
                signal performance_counter_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal performance_counter_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal performance_counter_control_slave_any_continuerequest :  STD_LOGIC;
                signal performance_counter_control_slave_arb_counter_enable :  STD_LOGIC;
                signal performance_counter_control_slave_arb_share_counter :  STD_LOGIC;
                signal performance_counter_control_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal performance_counter_control_slave_arb_share_set_values :  STD_LOGIC;
                signal performance_counter_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal performance_counter_control_slave_begins_xfer :  STD_LOGIC;
                signal performance_counter_control_slave_end_xfer :  STD_LOGIC;
                signal performance_counter_control_slave_firsttransfer :  STD_LOGIC;
                signal performance_counter_control_slave_grant_vector :  STD_LOGIC;
                signal performance_counter_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal performance_counter_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal performance_counter_control_slave_master_qreq_vector :  STD_LOGIC;
                signal performance_counter_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal performance_counter_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal performance_counter_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal performance_counter_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal performance_counter_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal performance_counter_control_slave_waits_for_read :  STD_LOGIC;
                signal performance_counter_control_slave_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_performance_counter_control_slave_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_performance_counter_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT performance_counter_control_slave_end_xfer;
    end if;

  end process;

  performance_counter_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_performance_counter_control_slave);
  --assign performance_counter_control_slave_readdata_from_sa = performance_counter_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  performance_counter_control_slave_readdata_from_sa <= performance_counter_control_slave_readdata;
  internal_cpuNios_data_master_requests_performance_counter_control_slave <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 6) & std_logic_vector'("000000")) = std_logic_vector'("100000000000100010000000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --registered rdv signal_name registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave assignment, which is an e_assign
  registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave <= cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register_in;
  --performance_counter_control_slave_arb_share_counter set values, which is an e_mux
  performance_counter_control_slave_arb_share_set_values <= std_logic'('1');
  --performance_counter_control_slave_non_bursting_master_requests mux, which is an e_mux
  performance_counter_control_slave_non_bursting_master_requests <= internal_cpuNios_data_master_requests_performance_counter_control_slave;
  --performance_counter_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  performance_counter_control_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --performance_counter_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  performance_counter_control_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(performance_counter_control_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(performance_counter_control_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(performance_counter_control_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(performance_counter_control_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --performance_counter_control_slave_allgrants all slave grants, which is an e_mux
  performance_counter_control_slave_allgrants <= performance_counter_control_slave_grant_vector;
  --performance_counter_control_slave_end_xfer assignment, which is an e_assign
  performance_counter_control_slave_end_xfer <= NOT ((performance_counter_control_slave_waits_for_read OR performance_counter_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_performance_counter_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_performance_counter_control_slave <= performance_counter_control_slave_end_xfer AND (((NOT performance_counter_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --performance_counter_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  performance_counter_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_performance_counter_control_slave AND performance_counter_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_performance_counter_control_slave AND NOT performance_counter_control_slave_non_bursting_master_requests));
  --performance_counter_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      performance_counter_control_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(performance_counter_control_slave_arb_counter_enable) = '1' then 
        performance_counter_control_slave_arb_share_counter <= performance_counter_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --performance_counter_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      performance_counter_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((performance_counter_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_performance_counter_control_slave)) OR ((end_xfer_arb_share_counter_term_performance_counter_control_slave AND NOT performance_counter_control_slave_non_bursting_master_requests)))) = '1' then 
        performance_counter_control_slave_slavearbiterlockenable <= performance_counter_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master performance_counter/control_slave arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= performance_counter_control_slave_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --performance_counter_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  performance_counter_control_slave_slavearbiterlockenable2 <= performance_counter_control_slave_arb_share_counter_next_value;
  --cpuNios/data_master performance_counter/control_slave arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= performance_counter_control_slave_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --performance_counter_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  performance_counter_control_slave_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_performance_counter_control_slave <= internal_cpuNios_data_master_requests_performance_counter_control_slave AND NOT ((((cpuNios_data_master_read AND (cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register))) OR (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write))));
  --cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register_in <= ((internal_cpuNios_data_master_granted_performance_counter_control_slave AND cpuNios_data_master_read) AND NOT performance_counter_control_slave_waits_for_read) AND NOT (cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register);
  --shift register p1 cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register) & A_ToStdLogicVector(cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register_in)));
  --cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register <= p1_cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register;
    end if;

  end process;

  --local readdatavalid cpuNios_data_master_read_data_valid_performance_counter_control_slave, which is an e_mux
  cpuNios_data_master_read_data_valid_performance_counter_control_slave <= cpuNios_data_master_read_data_valid_performance_counter_control_slave_shift_register;
  --performance_counter_control_slave_writedata mux, which is an e_mux
  performance_counter_control_slave_writedata <= cpuNios_data_master_writedata;
  --master is always granted when requested
  internal_cpuNios_data_master_granted_performance_counter_control_slave <= internal_cpuNios_data_master_qualified_request_performance_counter_control_slave;
  --cpuNios/data_master saved-grant performance_counter/control_slave, which is an e_assign
  cpuNios_data_master_saved_grant_performance_counter_control_slave <= internal_cpuNios_data_master_requests_performance_counter_control_slave;
  --allow new arb cycle for performance_counter/control_slave, which is an e_assign
  performance_counter_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  performance_counter_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  performance_counter_control_slave_master_qreq_vector <= std_logic'('1');
  performance_counter_control_slave_begintransfer <= performance_counter_control_slave_begins_xfer;
  --performance_counter_control_slave_reset_n assignment, which is an e_assign
  performance_counter_control_slave_reset_n <= reset_n;
  --performance_counter_control_slave_firsttransfer first transaction, which is an e_assign
  performance_counter_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(performance_counter_control_slave_begins_xfer) = '1'), performance_counter_control_slave_unreg_firsttransfer, performance_counter_control_slave_reg_firsttransfer);
  --performance_counter_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  performance_counter_control_slave_unreg_firsttransfer <= NOT ((performance_counter_control_slave_slavearbiterlockenable AND performance_counter_control_slave_any_continuerequest));
  --performance_counter_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      performance_counter_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(performance_counter_control_slave_begins_xfer) = '1' then 
        performance_counter_control_slave_reg_firsttransfer <= performance_counter_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --performance_counter_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  performance_counter_control_slave_beginbursttransfer_internal <= performance_counter_control_slave_begins_xfer;
  --performance_counter_control_slave_write assignment, which is an e_mux
  performance_counter_control_slave_write <= internal_cpuNios_data_master_granted_performance_counter_control_slave AND cpuNios_data_master_write;
  shifted_address_to_performance_counter_control_slave_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --performance_counter_control_slave_address mux, which is an e_mux
  performance_counter_control_slave_address <= A_EXT (A_SRL(shifted_address_to_performance_counter_control_slave_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --d1_performance_counter_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_performance_counter_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_performance_counter_control_slave_end_xfer <= performance_counter_control_slave_end_xfer;
    end if;

  end process;

  --performance_counter_control_slave_waits_for_read in a cycle, which is an e_mux
  performance_counter_control_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(performance_counter_control_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --performance_counter_control_slave_in_a_read_cycle assignment, which is an e_assign
  performance_counter_control_slave_in_a_read_cycle <= internal_cpuNios_data_master_granted_performance_counter_control_slave AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= performance_counter_control_slave_in_a_read_cycle;
  --performance_counter_control_slave_waits_for_write in a cycle, which is an e_mux
  performance_counter_control_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(performance_counter_control_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --performance_counter_control_slave_in_a_write_cycle assignment, which is an e_assign
  performance_counter_control_slave_in_a_write_cycle <= internal_cpuNios_data_master_granted_performance_counter_control_slave AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= performance_counter_control_slave_in_a_write_cycle;
  wait_for_performance_counter_control_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_performance_counter_control_slave <= internal_cpuNios_data_master_granted_performance_counter_control_slave;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_performance_counter_control_slave <= internal_cpuNios_data_master_qualified_request_performance_counter_control_slave;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_performance_counter_control_slave <= internal_cpuNios_data_master_requests_performance_counter_control_slave;
--synthesis translate_off
    --performance_counter/control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_sdram_s1_module;


architecture europa of rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_lcd_sgdma_descriptor_read_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_lcd_sgdma_descriptor_read_to_sdram_s1_module;


architecture europa of rdv_fifo_for_lcd_sgdma_descriptor_read_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_lcd_sgdma_m_read_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_lcd_sgdma_m_read_to_sdram_s1_module;


architecture europa of rdv_fifo_for_lcd_sgdma_m_read_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_tse_ddr_clock_bridge_m1_to_sdram_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_tse_ddr_clock_bridge_m1_to_sdram_s1_module;


architecture europa of rdv_fifo_for_tse_ddr_clock_bridge_m1_to_sdram_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sdram_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_ddr_clock_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_descriptor_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_descriptor_read_latency_counter : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_read : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_descriptor_write_write : IN STD_LOGIC;
                 signal lcd_sgdma_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_m_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal lcd_sgdma_m_read_latency_counter : IN STD_LOGIC;
                 signal lcd_sgdma_m_read_read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal sdram_s1_readdatavalid : IN STD_LOGIC;
                 signal sdram_s1_resetrequest_n : IN STD_LOGIC;
                 signal sdram_s1_waitrequest_n : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal tse_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal tse_ddr_clock_bridge_m1_latency_counter : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal cpu_ddr_clock_bridge_m1_granted_sdram_s1 : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_ddr_clock_bridge_m1_requests_sdram_s1 : OUT STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : OUT STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_granted_sdram_s1 : OUT STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal lcd_sgdma_descriptor_read_requests_sdram_s1 : OUT STD_LOGIC;
                 signal lcd_sgdma_descriptor_write_granted_sdram_s1 : OUT STD_LOGIC;
                 signal lcd_sgdma_descriptor_write_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal lcd_sgdma_descriptor_write_requests_sdram_s1 : OUT STD_LOGIC;
                 signal lcd_sgdma_m_read_granted_sdram_s1 : OUT STD_LOGIC;
                 signal lcd_sgdma_m_read_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal lcd_sgdma_m_read_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal lcd_sgdma_m_read_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal lcd_sgdma_m_read_requests_sdram_s1 : OUT STD_LOGIC;
                 signal sdram_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal sdram_s1_beginbursttransfer : OUT STD_LOGIC;
                 signal sdram_s1_burstcount : OUT STD_LOGIC;
                 signal sdram_s1_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal sdram_s1_read : OUT STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal sdram_s1_resetrequest_n_from_sa : OUT STD_LOGIC;
                 signal sdram_s1_waitrequest_n_from_sa : OUT STD_LOGIC;
                 signal sdram_s1_write : OUT STD_LOGIC;
                 signal sdram_s1_writedata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal tse_ddr_clock_bridge_m1_granted_sdram_s1 : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_requests_sdram_s1 : OUT STD_LOGIC
              );
end entity sdram_s1_arbitrator;


architecture europa of sdram_s1_arbitrator is
component rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_sdram_s1_module;

component rdv_fifo_for_lcd_sgdma_descriptor_read_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_lcd_sgdma_descriptor_read_to_sdram_s1_module;

component rdv_fifo_for_lcd_sgdma_m_read_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_lcd_sgdma_m_read_to_sdram_s1_module;

component rdv_fifo_for_tse_ddr_clock_bridge_m1_to_sdram_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_tse_ddr_clock_bridge_m1_to_sdram_s1_module;

                signal cpu_ddr_clock_bridge_m1_arbiterlock :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_byteenable_sdram_s1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_continuerequest :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_saved_grant_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_writedata_replicated :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sdram_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1 :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1 :  STD_LOGIC;
                signal internal_lcd_sgdma_descriptor_read_granted_sdram_s1 :  STD_LOGIC;
                signal internal_lcd_sgdma_descriptor_read_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_lcd_sgdma_descriptor_read_requests_sdram_s1 :  STD_LOGIC;
                signal internal_lcd_sgdma_descriptor_write_granted_sdram_s1 :  STD_LOGIC;
                signal internal_lcd_sgdma_descriptor_write_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_lcd_sgdma_descriptor_write_requests_sdram_s1 :  STD_LOGIC;
                signal internal_lcd_sgdma_m_read_granted_sdram_s1 :  STD_LOGIC;
                signal internal_lcd_sgdma_m_read_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_lcd_sgdma_m_read_requests_sdram_s1 :  STD_LOGIC;
                signal internal_sdram_s1_waitrequest_n_from_sa :  STD_LOGIC;
                signal internal_tse_ddr_clock_bridge_m1_granted_sdram_s1 :  STD_LOGIC;
                signal internal_tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 :  STD_LOGIC;
                signal internal_tse_ddr_clock_bridge_m1_requests_sdram_s1 :  STD_LOGIC;
                signal last_cycle_cpu_ddr_clock_bridge_m1_granted_slave_sdram_s1 :  STD_LOGIC;
                signal last_cycle_lcd_sgdma_descriptor_read_granted_slave_sdram_s1 :  STD_LOGIC;
                signal last_cycle_lcd_sgdma_descriptor_write_granted_slave_sdram_s1 :  STD_LOGIC;
                signal last_cycle_lcd_sgdma_m_read_granted_slave_sdram_s1 :  STD_LOGIC;
                signal last_cycle_tse_ddr_clock_bridge_m1_granted_slave_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_arbiterlock :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_arbiterlock2 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_continuerequest :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_saved_grant_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_arbiterlock :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_arbiterlock2 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_byteenable_sdram_s1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal lcd_sgdma_descriptor_write_continuerequest :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_saved_grant_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_writedata_replicated :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal lcd_sgdma_m_read_arbiterlock :  STD_LOGIC;
                signal lcd_sgdma_m_read_arbiterlock2 :  STD_LOGIC;
                signal lcd_sgdma_m_read_continuerequest :  STD_LOGIC;
                signal lcd_sgdma_m_read_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_m_read_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_m_read_saved_grant_sdram_s1 :  STD_LOGIC;
                signal module_input18 :  STD_LOGIC;
                signal module_input19 :  STD_LOGIC;
                signal module_input20 :  STD_LOGIC;
                signal module_input21 :  STD_LOGIC;
                signal module_input22 :  STD_LOGIC;
                signal module_input23 :  STD_LOGIC;
                signal module_input24 :  STD_LOGIC;
                signal module_input25 :  STD_LOGIC;
                signal module_input26 :  STD_LOGIC;
                signal module_input27 :  STD_LOGIC;
                signal module_input28 :  STD_LOGIC;
                signal module_input29 :  STD_LOGIC;
                signal sdram_s1_allgrants :  STD_LOGIC;
                signal sdram_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sdram_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sdram_s1_any_continuerequest :  STD_LOGIC;
                signal sdram_s1_arb_addend :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sdram_s1_arb_counter_enable :  STD_LOGIC;
                signal sdram_s1_arb_share_counter :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal sdram_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal sdram_s1_arb_share_set_values :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal sdram_s1_arb_winner :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sdram_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal sdram_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sdram_s1_begins_xfer :  STD_LOGIC;
                signal sdram_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal sdram_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sdram_s1_end_xfer :  STD_LOGIC;
                signal sdram_s1_firsttransfer :  STD_LOGIC;
                signal sdram_s1_grant_vector :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sdram_s1_in_a_read_cycle :  STD_LOGIC;
                signal sdram_s1_in_a_write_cycle :  STD_LOGIC;
                signal sdram_s1_master_qreq_vector :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sdram_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal sdram_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sdram_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal sdram_s1_reg_firsttransfer :  STD_LOGIC;
                signal sdram_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sdram_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sdram_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sdram_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sdram_s1_waits_for_read :  STD_LOGIC;
                signal sdram_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_sdram_s1_from_cpu_ddr_clock_bridge_m1 :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal shifted_address_to_sdram_s1_from_lcd_sgdma_descriptor_read :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_sdram_s1_from_lcd_sgdma_descriptor_write :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_sdram_s1_from_lcd_sgdma_m_read :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_sdram_s1_from_tse_ddr_clock_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal tse_ddr_clock_bridge_m1_arbiterlock :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_byteenable_sdram_s1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal tse_ddr_clock_bridge_m1_continuerequest :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_rdv_fifo_empty_sdram_s1 :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_rdv_fifo_output_from_sdram_s1 :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_saved_grant_sdram_s1 :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_writedata_replicated :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal wait_for_sdram_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sdram_s1_end_xfer;
    end if;

  end process;

  sdram_s1_begins_xfer <= NOT d1_reasons_to_wait AND (((((internal_cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 OR internal_lcd_sgdma_descriptor_read_qualified_request_sdram_s1) OR internal_lcd_sgdma_descriptor_write_qualified_request_sdram_s1) OR internal_lcd_sgdma_m_read_qualified_request_sdram_s1) OR internal_tse_ddr_clock_bridge_m1_qualified_request_sdram_s1));
  --assign sdram_s1_readdatavalid_from_sa = sdram_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_s1_readdatavalid_from_sa <= sdram_s1_readdatavalid;
  --assign sdram_s1_readdata_from_sa = sdram_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_s1_readdata_from_sa <= sdram_s1_readdata;
  internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1 <= to_std_logic(((Std_Logic_Vector'(A_ToStdLogicVector(cpu_ddr_clock_bridge_m1_address_to_slave(25)) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000000000000000000000000")))) AND ((cpu_ddr_clock_bridge_m1_read OR cpu_ddr_clock_bridge_m1_write));
  --assign sdram_s1_waitrequest_n_from_sa = sdram_s1_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_sdram_s1_waitrequest_n_from_sa <= sdram_s1_waitrequest_n;
  --sdram_s1_arb_share_counter set values, which is an e_mux
  sdram_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_read_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000001100100"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_write_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000001100100"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_m_read_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000110010"), A_WE_StdLogicVector((std_logic'((internal_tse_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_read_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000001100100"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_write_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000001100100"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_m_read_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000110010"), A_WE_StdLogicVector((std_logic'((internal_tse_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_read_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000001100100"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_write_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000001100100"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_m_read_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000110010"), A_WE_StdLogicVector((std_logic'((internal_tse_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_read_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000001100100"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_write_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000001100100"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_m_read_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000110010"), A_WE_StdLogicVector((std_logic'((internal_tse_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_read_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000001100100"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_write_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000001100100"), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_m_read_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000110010"), A_WE_StdLogicVector((std_logic'((internal_tse_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), std_logic_vector'("00000000000000000000000000000001")))))))))))))))))))))))))), 7);
  --sdram_s1_non_bursting_master_requests mux, which is an e_mux
  sdram_s1_non_bursting_master_requests <= (((((((((((((((((((((((internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1 OR internal_lcd_sgdma_descriptor_read_requests_sdram_s1) OR internal_lcd_sgdma_descriptor_write_requests_sdram_s1) OR internal_lcd_sgdma_m_read_requests_sdram_s1) OR internal_tse_ddr_clock_bridge_m1_requests_sdram_s1) OR internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1) OR internal_lcd_sgdma_descriptor_read_requests_sdram_s1) OR internal_lcd_sgdma_descriptor_write_requests_sdram_s1) OR internal_lcd_sgdma_m_read_requests_sdram_s1) OR internal_tse_ddr_clock_bridge_m1_requests_sdram_s1) OR internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1) OR internal_lcd_sgdma_descriptor_read_requests_sdram_s1) OR internal_lcd_sgdma_descriptor_write_requests_sdram_s1) OR internal_lcd_sgdma_m_read_requests_sdram_s1) OR internal_tse_ddr_clock_bridge_m1_requests_sdram_s1) OR internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1) OR internal_lcd_sgdma_descriptor_read_requests_sdram_s1) OR internal_lcd_sgdma_descriptor_write_requests_sdram_s1) OR internal_lcd_sgdma_m_read_requests_sdram_s1) OR internal_tse_ddr_clock_bridge_m1_requests_sdram_s1) OR internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1) OR internal_lcd_sgdma_descriptor_read_requests_sdram_s1) OR internal_lcd_sgdma_descriptor_write_requests_sdram_s1) OR internal_lcd_sgdma_m_read_requests_sdram_s1) OR internal_tse_ddr_clock_bridge_m1_requests_sdram_s1;
  --sdram_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sdram_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sdram_s1_arb_share_counter_next_value assignment, which is an e_assign
  sdram_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sdram_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000") & (sdram_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sdram_s1_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000") & (sdram_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 7);
  --sdram_s1_allgrants all slave grants, which is an e_mux
  sdram_s1_allgrants <= ((((((((((((((((((((((((or_reduce(sdram_s1_grant_vector)) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector))) OR (or_reduce(sdram_s1_grant_vector));
  --sdram_s1_end_xfer assignment, which is an e_assign
  sdram_s1_end_xfer <= NOT ((sdram_s1_waits_for_read OR sdram_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sdram_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sdram_s1 <= sdram_s1_end_xfer AND (((NOT sdram_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sdram_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sdram_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sdram_s1 AND sdram_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sdram_s1 AND NOT sdram_s1_non_bursting_master_requests));
  --sdram_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_arb_share_counter <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_arb_counter_enable) = '1' then 
        sdram_s1_arb_share_counter <= sdram_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sdram_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(sdram_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_sdram_s1)) OR ((end_xfer_arb_share_counter_term_sdram_s1 AND NOT sdram_s1_non_bursting_master_requests)))) = '1' then 
        sdram_s1_slavearbiterlockenable <= or_reduce(sdram_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu_ddr_clock_bridge/m1 sdram/s1 arbiterlock, which is an e_assign
  cpu_ddr_clock_bridge_m1_arbiterlock <= sdram_s1_slavearbiterlockenable AND cpu_ddr_clock_bridge_m1_continuerequest;
  --sdram_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sdram_s1_slavearbiterlockenable2 <= or_reduce(sdram_s1_arb_share_counter_next_value);
  --cpu_ddr_clock_bridge/m1 sdram/s1 arbiterlock2, which is an e_assign
  cpu_ddr_clock_bridge_m1_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND cpu_ddr_clock_bridge_m1_continuerequest;
  --lcd_sgdma/descriptor_read sdram/s1 arbiterlock, which is an e_assign
  lcd_sgdma_descriptor_read_arbiterlock <= sdram_s1_slavearbiterlockenable AND lcd_sgdma_descriptor_read_continuerequest;
  --lcd_sgdma/descriptor_read sdram/s1 arbiterlock2, which is an e_assign
  lcd_sgdma_descriptor_read_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND lcd_sgdma_descriptor_read_continuerequest;
  --lcd_sgdma/descriptor_read granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_lcd_sgdma_descriptor_read_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_lcd_sgdma_descriptor_read_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(lcd_sgdma_descriptor_read_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_s1_arbitration_holdoff_internal OR NOT internal_lcd_sgdma_descriptor_read_requests_sdram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_lcd_sgdma_descriptor_read_granted_slave_sdram_s1))))));
    end if;

  end process;

  --lcd_sgdma_descriptor_read_continuerequest continued request, which is an e_mux
  lcd_sgdma_descriptor_read_continuerequest <= ((((last_cycle_lcd_sgdma_descriptor_read_granted_slave_sdram_s1 AND internal_lcd_sgdma_descriptor_read_requests_sdram_s1)) OR ((last_cycle_lcd_sgdma_descriptor_read_granted_slave_sdram_s1 AND internal_lcd_sgdma_descriptor_read_requests_sdram_s1))) OR ((last_cycle_lcd_sgdma_descriptor_read_granted_slave_sdram_s1 AND internal_lcd_sgdma_descriptor_read_requests_sdram_s1))) OR ((last_cycle_lcd_sgdma_descriptor_read_granted_slave_sdram_s1 AND internal_lcd_sgdma_descriptor_read_requests_sdram_s1));
  --sdram_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  sdram_s1_any_continuerequest <= ((((((((((((((((((lcd_sgdma_descriptor_read_continuerequest OR lcd_sgdma_descriptor_write_continuerequest) OR lcd_sgdma_m_read_continuerequest) OR tse_ddr_clock_bridge_m1_continuerequest) OR cpu_ddr_clock_bridge_m1_continuerequest) OR lcd_sgdma_descriptor_write_continuerequest) OR lcd_sgdma_m_read_continuerequest) OR tse_ddr_clock_bridge_m1_continuerequest) OR cpu_ddr_clock_bridge_m1_continuerequest) OR lcd_sgdma_descriptor_read_continuerequest) OR lcd_sgdma_m_read_continuerequest) OR tse_ddr_clock_bridge_m1_continuerequest) OR cpu_ddr_clock_bridge_m1_continuerequest) OR lcd_sgdma_descriptor_read_continuerequest) OR lcd_sgdma_descriptor_write_continuerequest) OR tse_ddr_clock_bridge_m1_continuerequest) OR cpu_ddr_clock_bridge_m1_continuerequest) OR lcd_sgdma_descriptor_read_continuerequest) OR lcd_sgdma_descriptor_write_continuerequest) OR lcd_sgdma_m_read_continuerequest;
  --lcd_sgdma/descriptor_write sdram/s1 arbiterlock, which is an e_assign
  lcd_sgdma_descriptor_write_arbiterlock <= sdram_s1_slavearbiterlockenable AND lcd_sgdma_descriptor_write_continuerequest;
  --lcd_sgdma/descriptor_write sdram/s1 arbiterlock2, which is an e_assign
  lcd_sgdma_descriptor_write_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND lcd_sgdma_descriptor_write_continuerequest;
  --lcd_sgdma/descriptor_write granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_lcd_sgdma_descriptor_write_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_lcd_sgdma_descriptor_write_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(lcd_sgdma_descriptor_write_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_s1_arbitration_holdoff_internal OR NOT internal_lcd_sgdma_descriptor_write_requests_sdram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_lcd_sgdma_descriptor_write_granted_slave_sdram_s1))))));
    end if;

  end process;

  --lcd_sgdma_descriptor_write_continuerequest continued request, which is an e_mux
  lcd_sgdma_descriptor_write_continuerequest <= ((((last_cycle_lcd_sgdma_descriptor_write_granted_slave_sdram_s1 AND internal_lcd_sgdma_descriptor_write_requests_sdram_s1)) OR ((last_cycle_lcd_sgdma_descriptor_write_granted_slave_sdram_s1 AND internal_lcd_sgdma_descriptor_write_requests_sdram_s1))) OR ((last_cycle_lcd_sgdma_descriptor_write_granted_slave_sdram_s1 AND internal_lcd_sgdma_descriptor_write_requests_sdram_s1))) OR ((last_cycle_lcd_sgdma_descriptor_write_granted_slave_sdram_s1 AND internal_lcd_sgdma_descriptor_write_requests_sdram_s1));
  --lcd_sgdma/m_read sdram/s1 arbiterlock, which is an e_assign
  lcd_sgdma_m_read_arbiterlock <= sdram_s1_slavearbiterlockenable AND lcd_sgdma_m_read_continuerequest;
  --lcd_sgdma/m_read sdram/s1 arbiterlock2, which is an e_assign
  lcd_sgdma_m_read_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND lcd_sgdma_m_read_continuerequest;
  --lcd_sgdma/m_read granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_lcd_sgdma_m_read_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_lcd_sgdma_m_read_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(lcd_sgdma_m_read_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_s1_arbitration_holdoff_internal OR NOT internal_lcd_sgdma_m_read_requests_sdram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_lcd_sgdma_m_read_granted_slave_sdram_s1))))));
    end if;

  end process;

  --lcd_sgdma_m_read_continuerequest continued request, which is an e_mux
  lcd_sgdma_m_read_continuerequest <= ((((last_cycle_lcd_sgdma_m_read_granted_slave_sdram_s1 AND internal_lcd_sgdma_m_read_requests_sdram_s1)) OR ((last_cycle_lcd_sgdma_m_read_granted_slave_sdram_s1 AND internal_lcd_sgdma_m_read_requests_sdram_s1))) OR ((last_cycle_lcd_sgdma_m_read_granted_slave_sdram_s1 AND internal_lcd_sgdma_m_read_requests_sdram_s1))) OR ((last_cycle_lcd_sgdma_m_read_granted_slave_sdram_s1 AND internal_lcd_sgdma_m_read_requests_sdram_s1));
  --tse_ddr_clock_bridge/m1 sdram/s1 arbiterlock, which is an e_assign
  tse_ddr_clock_bridge_m1_arbiterlock <= sdram_s1_slavearbiterlockenable AND tse_ddr_clock_bridge_m1_continuerequest;
  --tse_ddr_clock_bridge/m1 sdram/s1 arbiterlock2, which is an e_assign
  tse_ddr_clock_bridge_m1_arbiterlock2 <= sdram_s1_slavearbiterlockenable2 AND tse_ddr_clock_bridge_m1_continuerequest;
  --tse_ddr_clock_bridge/m1 granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_tse_ddr_clock_bridge_m1_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_tse_ddr_clock_bridge_m1_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(tse_ddr_clock_bridge_m1_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_s1_arbitration_holdoff_internal OR NOT internal_tse_ddr_clock_bridge_m1_requests_sdram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_tse_ddr_clock_bridge_m1_granted_slave_sdram_s1))))));
    end if;

  end process;

  --tse_ddr_clock_bridge_m1_continuerequest continued request, which is an e_mux
  tse_ddr_clock_bridge_m1_continuerequest <= ((((last_cycle_tse_ddr_clock_bridge_m1_granted_slave_sdram_s1 AND internal_tse_ddr_clock_bridge_m1_requests_sdram_s1)) OR ((last_cycle_tse_ddr_clock_bridge_m1_granted_slave_sdram_s1 AND internal_tse_ddr_clock_bridge_m1_requests_sdram_s1))) OR ((last_cycle_tse_ddr_clock_bridge_m1_granted_slave_sdram_s1 AND internal_tse_ddr_clock_bridge_m1_requests_sdram_s1))) OR ((last_cycle_tse_ddr_clock_bridge_m1_granted_slave_sdram_s1 AND internal_tse_ddr_clock_bridge_m1_requests_sdram_s1));
  internal_cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 <= internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1 AND NOT (((((((cpu_ddr_clock_bridge_m1_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_m1_latency_counter)))))))))) OR lcd_sgdma_descriptor_read_arbiterlock) OR lcd_sgdma_descriptor_write_arbiterlock) OR lcd_sgdma_m_read_arbiterlock) OR tse_ddr_clock_bridge_m1_arbiterlock));
  --unique name for sdram_s1_move_on_to_next_transaction, which is an e_assign
  sdram_s1_move_on_to_next_transaction <= sdram_s1_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_sdram_s1 : rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_sdram_s1_module
    port map(
      data_out => cpu_ddr_clock_bridge_m1_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => cpu_ddr_clock_bridge_m1_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input18,
      clk => clk,
      data_in => internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input19,
      write => module_input20
    );

  module_input18 <= std_logic'('0');
  module_input19 <= std_logic'('0');
  module_input20 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register <= NOT cpu_ddr_clock_bridge_m1_rdv_fifo_empty_sdram_s1;
  --local readdatavalid cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1, which is an e_mux
  cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND cpu_ddr_clock_bridge_m1_rdv_fifo_output_from_sdram_s1)) AND NOT cpu_ddr_clock_bridge_m1_rdv_fifo_empty_sdram_s1;
  --replicate narrow data for wide slave
  cpu_ddr_clock_bridge_m1_writedata_replicated <= cpu_ddr_clock_bridge_m1_writedata & cpu_ddr_clock_bridge_m1_writedata;
  --sdram_s1_writedata mux, which is an e_mux
  sdram_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), cpu_ddr_clock_bridge_m1_writedata_replicated, A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_write_granted_sdram_s1)) = '1'), lcd_sgdma_descriptor_write_writedata_replicated, tse_ddr_clock_bridge_m1_writedata_replicated));
  internal_lcd_sgdma_descriptor_read_requests_sdram_s1 <= ((to_std_logic(((Std_Logic_Vector'(lcd_sgdma_descriptor_read_address_to_slave(31 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (lcd_sgdma_descriptor_read_read))) AND lcd_sgdma_descriptor_read_read;
  --cpu_ddr_clock_bridge/m1 granted sdram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_ddr_clock_bridge_m1_granted_slave_sdram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_ddr_clock_bridge_m1_granted_slave_sdram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_ddr_clock_bridge_m1_saved_grant_sdram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_s1_arbitration_holdoff_internal OR NOT internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_ddr_clock_bridge_m1_granted_slave_sdram_s1))))));
    end if;

  end process;

  --cpu_ddr_clock_bridge_m1_continuerequest continued request, which is an e_mux
  cpu_ddr_clock_bridge_m1_continuerequest <= ((((last_cycle_cpu_ddr_clock_bridge_m1_granted_slave_sdram_s1 AND internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1)) OR ((last_cycle_cpu_ddr_clock_bridge_m1_granted_slave_sdram_s1 AND internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1))) OR ((last_cycle_cpu_ddr_clock_bridge_m1_granted_slave_sdram_s1 AND internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1))) OR ((last_cycle_cpu_ddr_clock_bridge_m1_granted_slave_sdram_s1 AND internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1));
  internal_lcd_sgdma_descriptor_read_qualified_request_sdram_s1 <= internal_lcd_sgdma_descriptor_read_requests_sdram_s1 AND NOT (((((((lcd_sgdma_descriptor_read_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_sgdma_descriptor_read_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_sgdma_descriptor_read_latency_counter)))))))))) OR cpu_ddr_clock_bridge_m1_arbiterlock) OR lcd_sgdma_descriptor_write_arbiterlock) OR lcd_sgdma_m_read_arbiterlock) OR tse_ddr_clock_bridge_m1_arbiterlock));
  --rdv_fifo_for_lcd_sgdma_descriptor_read_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_lcd_sgdma_descriptor_read_to_sdram_s1 : rdv_fifo_for_lcd_sgdma_descriptor_read_to_sdram_s1_module
    port map(
      data_out => lcd_sgdma_descriptor_read_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => lcd_sgdma_descriptor_read_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input21,
      clk => clk,
      data_in => internal_lcd_sgdma_descriptor_read_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input22,
      write => module_input23
    );

  module_input21 <= std_logic'('0');
  module_input22 <= std_logic'('0');
  module_input23 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  lcd_sgdma_descriptor_read_read_data_valid_sdram_s1_shift_register <= NOT lcd_sgdma_descriptor_read_rdv_fifo_empty_sdram_s1;
  --local readdatavalid lcd_sgdma_descriptor_read_read_data_valid_sdram_s1, which is an e_mux
  lcd_sgdma_descriptor_read_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND lcd_sgdma_descriptor_read_rdv_fifo_output_from_sdram_s1)) AND NOT lcd_sgdma_descriptor_read_rdv_fifo_empty_sdram_s1;
  internal_lcd_sgdma_descriptor_write_requests_sdram_s1 <= ((to_std_logic(((Std_Logic_Vector'(lcd_sgdma_descriptor_write_address_to_slave(31 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (lcd_sgdma_descriptor_write_write))) AND lcd_sgdma_descriptor_write_write;
  internal_lcd_sgdma_descriptor_write_qualified_request_sdram_s1 <= internal_lcd_sgdma_descriptor_write_requests_sdram_s1 AND NOT ((((cpu_ddr_clock_bridge_m1_arbiterlock OR lcd_sgdma_descriptor_read_arbiterlock) OR lcd_sgdma_m_read_arbiterlock) OR tse_ddr_clock_bridge_m1_arbiterlock));
  --replicate narrow data for wide slave
  lcd_sgdma_descriptor_write_writedata_replicated <= lcd_sgdma_descriptor_write_writedata & lcd_sgdma_descriptor_write_writedata;
  internal_lcd_sgdma_m_read_requests_sdram_s1 <= ((to_std_logic(((Std_Logic_Vector'(lcd_sgdma_m_read_address_to_slave(31 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (lcd_sgdma_m_read_read))) AND lcd_sgdma_m_read_read;
  internal_lcd_sgdma_m_read_qualified_request_sdram_s1 <= internal_lcd_sgdma_m_read_requests_sdram_s1 AND NOT (((((((lcd_sgdma_m_read_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_sgdma_m_read_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_sgdma_m_read_latency_counter)))))))))) OR cpu_ddr_clock_bridge_m1_arbiterlock) OR lcd_sgdma_descriptor_read_arbiterlock) OR lcd_sgdma_descriptor_write_arbiterlock) OR tse_ddr_clock_bridge_m1_arbiterlock));
  --rdv_fifo_for_lcd_sgdma_m_read_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_lcd_sgdma_m_read_to_sdram_s1 : rdv_fifo_for_lcd_sgdma_m_read_to_sdram_s1_module
    port map(
      data_out => lcd_sgdma_m_read_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => lcd_sgdma_m_read_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input24,
      clk => clk,
      data_in => internal_lcd_sgdma_m_read_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input25,
      write => module_input26
    );

  module_input24 <= std_logic'('0');
  module_input25 <= std_logic'('0');
  module_input26 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  lcd_sgdma_m_read_read_data_valid_sdram_s1_shift_register <= NOT lcd_sgdma_m_read_rdv_fifo_empty_sdram_s1;
  --local readdatavalid lcd_sgdma_m_read_read_data_valid_sdram_s1, which is an e_mux
  lcd_sgdma_m_read_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND lcd_sgdma_m_read_rdv_fifo_output_from_sdram_s1)) AND NOT lcd_sgdma_m_read_rdv_fifo_empty_sdram_s1;
  internal_tse_ddr_clock_bridge_m1_requests_sdram_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((tse_ddr_clock_bridge_m1_read OR tse_ddr_clock_bridge_m1_write)))))));
  internal_tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 <= internal_tse_ddr_clock_bridge_m1_requests_sdram_s1 AND NOT (((((((tse_ddr_clock_bridge_m1_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_ddr_clock_bridge_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_ddr_clock_bridge_m1_latency_counter)))))))))) OR cpu_ddr_clock_bridge_m1_arbiterlock) OR lcd_sgdma_descriptor_read_arbiterlock) OR lcd_sgdma_descriptor_write_arbiterlock) OR lcd_sgdma_m_read_arbiterlock));
  --rdv_fifo_for_tse_ddr_clock_bridge_m1_to_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_tse_ddr_clock_bridge_m1_to_sdram_s1 : rdv_fifo_for_tse_ddr_clock_bridge_m1_to_sdram_s1_module
    port map(
      data_out => tse_ddr_clock_bridge_m1_rdv_fifo_output_from_sdram_s1,
      empty => open,
      fifo_contains_ones_n => tse_ddr_clock_bridge_m1_rdv_fifo_empty_sdram_s1,
      full => open,
      clear_fifo => module_input27,
      clk => clk,
      data_in => internal_tse_ddr_clock_bridge_m1_granted_sdram_s1,
      read => sdram_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input28,
      write => module_input29
    );

  module_input27 <= std_logic'('0');
  module_input28 <= std_logic'('0');
  module_input29 <= in_a_read_cycle AND NOT sdram_s1_waits_for_read;

  tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register <= NOT tse_ddr_clock_bridge_m1_rdv_fifo_empty_sdram_s1;
  --local readdatavalid tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1, which is an e_mux
  tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1 <= ((sdram_s1_readdatavalid_from_sa AND tse_ddr_clock_bridge_m1_rdv_fifo_output_from_sdram_s1)) AND NOT tse_ddr_clock_bridge_m1_rdv_fifo_empty_sdram_s1;
  --replicate narrow data for wide slave
  tse_ddr_clock_bridge_m1_writedata_replicated <= tse_ddr_clock_bridge_m1_writedata & tse_ddr_clock_bridge_m1_writedata;
  --allow new arb cycle for sdram/s1, which is an e_assign
  sdram_s1_allow_new_arb_cycle <= (((NOT cpu_ddr_clock_bridge_m1_arbiterlock AND NOT lcd_sgdma_descriptor_read_arbiterlock) AND NOT lcd_sgdma_descriptor_write_arbiterlock) AND NOT lcd_sgdma_m_read_arbiterlock) AND NOT tse_ddr_clock_bridge_m1_arbiterlock;
  --tse_ddr_clock_bridge/m1 assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(0) <= internal_tse_ddr_clock_bridge_m1_qualified_request_sdram_s1;
  --tse_ddr_clock_bridge/m1 grant sdram/s1, which is an e_assign
  internal_tse_ddr_clock_bridge_m1_granted_sdram_s1 <= sdram_s1_grant_vector(0);
  --tse_ddr_clock_bridge/m1 saved-grant sdram/s1, which is an e_assign
  tse_ddr_clock_bridge_m1_saved_grant_sdram_s1 <= sdram_s1_arb_winner(0) AND internal_tse_ddr_clock_bridge_m1_requests_sdram_s1;
  --lcd_sgdma/m_read assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(1) <= internal_lcd_sgdma_m_read_qualified_request_sdram_s1;
  --lcd_sgdma/m_read grant sdram/s1, which is an e_assign
  internal_lcd_sgdma_m_read_granted_sdram_s1 <= sdram_s1_grant_vector(1);
  --lcd_sgdma/m_read saved-grant sdram/s1, which is an e_assign
  lcd_sgdma_m_read_saved_grant_sdram_s1 <= sdram_s1_arb_winner(1) AND internal_lcd_sgdma_m_read_requests_sdram_s1;
  --lcd_sgdma/descriptor_write assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(2) <= internal_lcd_sgdma_descriptor_write_qualified_request_sdram_s1;
  --lcd_sgdma/descriptor_write grant sdram/s1, which is an e_assign
  internal_lcd_sgdma_descriptor_write_granted_sdram_s1 <= sdram_s1_grant_vector(2);
  --lcd_sgdma/descriptor_write saved-grant sdram/s1, which is an e_assign
  lcd_sgdma_descriptor_write_saved_grant_sdram_s1 <= sdram_s1_arb_winner(2) AND internal_lcd_sgdma_descriptor_write_requests_sdram_s1;
  --lcd_sgdma/descriptor_read assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(3) <= internal_lcd_sgdma_descriptor_read_qualified_request_sdram_s1;
  --lcd_sgdma/descriptor_read grant sdram/s1, which is an e_assign
  internal_lcd_sgdma_descriptor_read_granted_sdram_s1 <= sdram_s1_grant_vector(3);
  --lcd_sgdma/descriptor_read saved-grant sdram/s1, which is an e_assign
  lcd_sgdma_descriptor_read_saved_grant_sdram_s1 <= sdram_s1_arb_winner(3) AND internal_lcd_sgdma_descriptor_read_requests_sdram_s1;
  --cpu_ddr_clock_bridge/m1 assignment into master qualified-requests vector for sdram/s1, which is an e_assign
  sdram_s1_master_qreq_vector(4) <= internal_cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1;
  --cpu_ddr_clock_bridge/m1 grant sdram/s1, which is an e_assign
  internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1 <= sdram_s1_grant_vector(4);
  --cpu_ddr_clock_bridge/m1 saved-grant sdram/s1, which is an e_assign
  cpu_ddr_clock_bridge_m1_saved_grant_sdram_s1 <= sdram_s1_arb_winner(4) AND internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1;
  --sdram/s1 chosen-master double-vector, which is an e_assign
  sdram_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((sdram_s1_master_qreq_vector & sdram_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT sdram_s1_master_qreq_vector & NOT sdram_s1_master_qreq_vector))) + (std_logic_vector'("000000") & (sdram_s1_arb_addend))))), 10);
  --stable onehot encoding of arb winner
  sdram_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((sdram_s1_allow_new_arb_cycle AND or_reduce(sdram_s1_grant_vector)))) = '1'), sdram_s1_grant_vector, sdram_s1_saved_chosen_master_vector);
  --saved sdram_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_saved_chosen_master_vector <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_allow_new_arb_cycle) = '1' then 
        sdram_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(sdram_s1_grant_vector)) = '1'), sdram_s1_grant_vector, sdram_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  sdram_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(4) OR sdram_s1_chosen_master_double_vector(9)))) & A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(3) OR sdram_s1_chosen_master_double_vector(8)))) & A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(2) OR sdram_s1_chosen_master_double_vector(7)))) & A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(1) OR sdram_s1_chosen_master_double_vector(6)))) & A_ToStdLogicVector(((sdram_s1_chosen_master_double_vector(0) OR sdram_s1_chosen_master_double_vector(5)))));
  --sdram/s1 chosen master rotated left, which is an e_assign
  sdram_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(sdram_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00000")), (std_logic_vector'("000000000000000000000000000") & ((A_SLL(sdram_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 5);
  --sdram/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_arb_addend <= std_logic_vector'("00001");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(sdram_s1_grant_vector)) = '1' then 
        sdram_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(sdram_s1_end_xfer) = '1'), sdram_s1_chosen_master_rot_left, sdram_s1_grant_vector);
      end if;
    end if;

  end process;

  --assign sdram_s1_resetrequest_n_from_sa = sdram_s1_resetrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_s1_resetrequest_n_from_sa <= sdram_s1_resetrequest_n;
  --sdram_s1_firsttransfer first transaction, which is an e_assign
  sdram_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sdram_s1_begins_xfer) = '1'), sdram_s1_unreg_firsttransfer, sdram_s1_reg_firsttransfer);
  --sdram_s1_unreg_firsttransfer first transaction, which is an e_assign
  sdram_s1_unreg_firsttransfer <= NOT ((sdram_s1_slavearbiterlockenable AND sdram_s1_any_continuerequest));
  --sdram_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_s1_begins_xfer) = '1' then 
        sdram_s1_reg_firsttransfer <= sdram_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sdram_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sdram_s1_beginbursttransfer_internal <= sdram_s1_begins_xfer;
  --sdram/s1 begin burst transfer to slave, which is an e_assign
  sdram_s1_beginbursttransfer <= sdram_s1_beginbursttransfer_internal;
  --sdram_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  sdram_s1_arbitration_holdoff_internal <= sdram_s1_begins_xfer AND sdram_s1_firsttransfer;
  --sdram_s1_read assignment, which is an e_mux
  sdram_s1_read <= ((((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1 AND cpu_ddr_clock_bridge_m1_read)) OR ((internal_lcd_sgdma_descriptor_read_granted_sdram_s1 AND lcd_sgdma_descriptor_read_read))) OR ((internal_lcd_sgdma_m_read_granted_sdram_s1 AND lcd_sgdma_m_read_read))) OR ((internal_tse_ddr_clock_bridge_m1_granted_sdram_s1 AND tse_ddr_clock_bridge_m1_read));
  --sdram_s1_write assignment, which is an e_mux
  sdram_s1_write <= (((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1 AND cpu_ddr_clock_bridge_m1_write)) OR ((internal_lcd_sgdma_descriptor_write_granted_sdram_s1 AND lcd_sgdma_descriptor_write_write))) OR ((internal_tse_ddr_clock_bridge_m1_granted_sdram_s1 AND tse_ddr_clock_bridge_m1_write));
  shifted_address_to_sdram_s1_from_cpu_ddr_clock_bridge_m1 <= cpu_ddr_clock_bridge_m1_address_to_slave;
  --sdram_s1_address mux, which is an e_mux
  sdram_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), (std_logic_vector'("000000") & ((A_SRL(shifted_address_to_sdram_s1_from_cpu_ddr_clock_bridge_m1,std_logic_vector'("00000000000000000000000000000011"))))), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_read_granted_sdram_s1)) = '1'), (A_SRL(shifted_address_to_sdram_s1_from_lcd_sgdma_descriptor_read,std_logic_vector'("00000000000000000000000000000011"))), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_write_granted_sdram_s1)) = '1'), (A_SRL(shifted_address_to_sdram_s1_from_lcd_sgdma_descriptor_write,std_logic_vector'("00000000000000000000000000000011"))), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_m_read_granted_sdram_s1)) = '1'), (A_SRL(shifted_address_to_sdram_s1_from_lcd_sgdma_m_read,std_logic_vector'("00000000000000000000000000000011"))), (std_logic_vector'("0000000") & ((A_SRL(shifted_address_to_sdram_s1_from_tse_ddr_clock_bridge_m1,std_logic_vector'("00000000000000000000000000000011"))))))))), 22);
  shifted_address_to_sdram_s1_from_lcd_sgdma_descriptor_read <= lcd_sgdma_descriptor_read_address_to_slave;
  shifted_address_to_sdram_s1_from_lcd_sgdma_descriptor_write <= lcd_sgdma_descriptor_write_address_to_slave;
  shifted_address_to_sdram_s1_from_lcd_sgdma_m_read <= lcd_sgdma_m_read_address_to_slave;
  shifted_address_to_sdram_s1_from_tse_ddr_clock_bridge_m1 <= tse_ddr_clock_bridge_m1_address_to_slave;
  --d1_sdram_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sdram_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sdram_s1_end_xfer <= sdram_s1_end_xfer;
    end if;

  end process;

  --sdram_s1_waits_for_read in a cycle, which is an e_mux
  sdram_s1_waits_for_read <= sdram_s1_in_a_read_cycle AND NOT internal_sdram_s1_waitrequest_n_from_sa;
  --sdram_s1_in_a_read_cycle assignment, which is an e_assign
  sdram_s1_in_a_read_cycle <= ((((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1 AND cpu_ddr_clock_bridge_m1_read)) OR ((internal_lcd_sgdma_descriptor_read_granted_sdram_s1 AND lcd_sgdma_descriptor_read_read))) OR ((internal_lcd_sgdma_m_read_granted_sdram_s1 AND lcd_sgdma_m_read_read))) OR ((internal_tse_ddr_clock_bridge_m1_granted_sdram_s1 AND tse_ddr_clock_bridge_m1_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sdram_s1_in_a_read_cycle;
  --sdram_s1_waits_for_write in a cycle, which is an e_mux
  sdram_s1_waits_for_write <= sdram_s1_in_a_write_cycle AND NOT internal_sdram_s1_waitrequest_n_from_sa;
  --sdram_s1_in_a_write_cycle assignment, which is an e_assign
  sdram_s1_in_a_write_cycle <= (((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1 AND cpu_ddr_clock_bridge_m1_write)) OR ((internal_lcd_sgdma_descriptor_write_granted_sdram_s1 AND lcd_sgdma_descriptor_write_write))) OR ((internal_tse_ddr_clock_bridge_m1_granted_sdram_s1 AND tse_ddr_clock_bridge_m1_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sdram_s1_in_a_write_cycle;
  wait_for_sdram_s1_counter <= std_logic'('0');
  --sdram_s1_byteenable byte enable port mux, which is an e_mux
  sdram_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000") & (cpu_ddr_clock_bridge_m1_byteenable_sdram_s1)), A_WE_StdLogicVector((std_logic'((internal_lcd_sgdma_descriptor_write_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000") & (lcd_sgdma_descriptor_write_byteenable_sdram_s1)), A_WE_StdLogicVector((std_logic'((internal_tse_ddr_clock_bridge_m1_granted_sdram_s1)) = '1'), (std_logic_vector'("000000000000000000000000") & (tse_ddr_clock_bridge_m1_byteenable_sdram_s1)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))))), 8);
  --byte_enable_mux for cpu_ddr_clock_bridge/m1 and sdram/s1, which is an e_mux
  cpu_ddr_clock_bridge_m1_byteenable_sdram_s1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_m1_address_to_slave(2)))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000") & (cpu_ddr_clock_bridge_m1_byteenable)), (cpu_ddr_clock_bridge_m1_byteenable & std_logic_vector'("0000")));
  --byte_enable_mux for lcd_sgdma/descriptor_write and sdram/s1, which is an e_mux
  lcd_sgdma_descriptor_write_byteenable_sdram_s1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(lcd_sgdma_descriptor_write_address_to_slave(2)))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000") & (A_REP(std_logic'('1'), 4))), (A_REP(std_logic'('1'), 4) & std_logic_vector'("0000")));
  --byte_enable_mux for tse_ddr_clock_bridge/m1 and sdram/s1, which is an e_mux
  tse_ddr_clock_bridge_m1_byteenable_sdram_s1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_ddr_clock_bridge_m1_address_to_slave(2)))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000") & (tse_ddr_clock_bridge_m1_byteenable)), (tse_ddr_clock_bridge_m1_byteenable & std_logic_vector'("0000")));
  --burstcount mux, which is an e_mux
  sdram_s1_burstcount <= std_logic'('1');
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_granted_sdram_s1 <= internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 <= internal_cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  cpu_ddr_clock_bridge_m1_requests_sdram_s1 <= internal_cpu_ddr_clock_bridge_m1_requests_sdram_s1;
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_read_granted_sdram_s1 <= internal_lcd_sgdma_descriptor_read_granted_sdram_s1;
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_read_qualified_request_sdram_s1 <= internal_lcd_sgdma_descriptor_read_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_read_requests_sdram_s1 <= internal_lcd_sgdma_descriptor_read_requests_sdram_s1;
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_write_granted_sdram_s1 <= internal_lcd_sgdma_descriptor_write_granted_sdram_s1;
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_write_qualified_request_sdram_s1 <= internal_lcd_sgdma_descriptor_write_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  lcd_sgdma_descriptor_write_requests_sdram_s1 <= internal_lcd_sgdma_descriptor_write_requests_sdram_s1;
  --vhdl renameroo for output signals
  lcd_sgdma_m_read_granted_sdram_s1 <= internal_lcd_sgdma_m_read_granted_sdram_s1;
  --vhdl renameroo for output signals
  lcd_sgdma_m_read_qualified_request_sdram_s1 <= internal_lcd_sgdma_m_read_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  lcd_sgdma_m_read_requests_sdram_s1 <= internal_lcd_sgdma_m_read_requests_sdram_s1;
  --vhdl renameroo for output signals
  sdram_s1_waitrequest_n_from_sa <= internal_sdram_s1_waitrequest_n_from_sa;
  --vhdl renameroo for output signals
  tse_ddr_clock_bridge_m1_granted_sdram_s1 <= internal_tse_ddr_clock_bridge_m1_granted_sdram_s1;
  --vhdl renameroo for output signals
  tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 <= internal_tse_ddr_clock_bridge_m1_qualified_request_sdram_s1;
  --vhdl renameroo for output signals
  tse_ddr_clock_bridge_m1_requests_sdram_s1 <= internal_tse_ddr_clock_bridge_m1_requests_sdram_s1;
--synthesis translate_off
    --sdram/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line34 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_ddr_clock_bridge_m1_granted_sdram_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_lcd_sgdma_descriptor_read_granted_sdram_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(internal_lcd_sgdma_descriptor_write_granted_sdram_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(internal_lcd_sgdma_m_read_granted_sdram_s1)))))) + (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(internal_tse_ddr_clock_bridge_m1_granted_sdram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line34, now);
          write(write_line34, string'(": "));
          write(write_line34, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line34.all);
          deallocate (write_line34);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line35 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_ddr_clock_bridge_m1_saved_grant_sdram_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(lcd_sgdma_descriptor_read_saved_grant_sdram_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(lcd_sgdma_descriptor_write_saved_grant_sdram_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(lcd_sgdma_m_read_saved_grant_sdram_s1)))))) + (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(tse_ddr_clock_bridge_m1_saved_grant_sdram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line35, now);
          write(write_line35, string'(": "));
          write(write_line35, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line35.all);
          deallocate (write_line35);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity processador_reset_clk50Mhz_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity processador_reset_clk50Mhz_domain_synch_module;


architecture europa of processador_reset_clk50Mhz_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sgdma_rx_csr_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_csr_irq : IN STD_LOGIC;
                 signal sgdma_rx_csr_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal cpuNios_data_master_granted_sgdma_rx_csr : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_sgdma_rx_csr : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_sgdma_rx_csr : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_sgdma_rx_csr : OUT STD_LOGIC;
                 signal d1_sgdma_rx_csr_end_xfer : OUT STD_LOGIC;
                 signal sgdma_rx_csr_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal sgdma_rx_csr_chipselect : OUT STD_LOGIC;
                 signal sgdma_rx_csr_irq_from_sa : OUT STD_LOGIC;
                 signal sgdma_rx_csr_read : OUT STD_LOGIC;
                 signal sgdma_rx_csr_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_csr_reset_n : OUT STD_LOGIC;
                 signal sgdma_rx_csr_write : OUT STD_LOGIC;
                 signal sgdma_rx_csr_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity sgdma_rx_csr_arbitrator;


architecture europa of sgdma_rx_csr_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_sgdma_rx_csr :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sgdma_rx_csr :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_sgdma_rx_csr :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_sgdma_rx_csr :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_sgdma_rx_csr :  STD_LOGIC;
                signal sgdma_rx_csr_allgrants :  STD_LOGIC;
                signal sgdma_rx_csr_allow_new_arb_cycle :  STD_LOGIC;
                signal sgdma_rx_csr_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sgdma_rx_csr_any_continuerequest :  STD_LOGIC;
                signal sgdma_rx_csr_arb_counter_enable :  STD_LOGIC;
                signal sgdma_rx_csr_arb_share_counter :  STD_LOGIC;
                signal sgdma_rx_csr_arb_share_counter_next_value :  STD_LOGIC;
                signal sgdma_rx_csr_arb_share_set_values :  STD_LOGIC;
                signal sgdma_rx_csr_beginbursttransfer_internal :  STD_LOGIC;
                signal sgdma_rx_csr_begins_xfer :  STD_LOGIC;
                signal sgdma_rx_csr_end_xfer :  STD_LOGIC;
                signal sgdma_rx_csr_firsttransfer :  STD_LOGIC;
                signal sgdma_rx_csr_grant_vector :  STD_LOGIC;
                signal sgdma_rx_csr_in_a_read_cycle :  STD_LOGIC;
                signal sgdma_rx_csr_in_a_write_cycle :  STD_LOGIC;
                signal sgdma_rx_csr_master_qreq_vector :  STD_LOGIC;
                signal sgdma_rx_csr_non_bursting_master_requests :  STD_LOGIC;
                signal sgdma_rx_csr_reg_firsttransfer :  STD_LOGIC;
                signal sgdma_rx_csr_slavearbiterlockenable :  STD_LOGIC;
                signal sgdma_rx_csr_slavearbiterlockenable2 :  STD_LOGIC;
                signal sgdma_rx_csr_unreg_firsttransfer :  STD_LOGIC;
                signal sgdma_rx_csr_waits_for_read :  STD_LOGIC;
                signal sgdma_rx_csr_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_sgdma_rx_csr_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_sgdma_rx_csr_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sgdma_rx_csr_end_xfer;
    end if;

  end process;

  sgdma_rx_csr_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_sgdma_rx_csr);
  --assign sgdma_rx_csr_readdata_from_sa = sgdma_rx_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sgdma_rx_csr_readdata_from_sa <= sgdma_rx_csr_readdata;
  internal_cpuNios_data_master_requests_sgdma_rx_csr <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 6) & std_logic_vector'("000000")) = std_logic_vector'("100000000000100100100000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --sgdma_rx_csr_arb_share_counter set values, which is an e_mux
  sgdma_rx_csr_arb_share_set_values <= std_logic'('1');
  --sgdma_rx_csr_non_bursting_master_requests mux, which is an e_mux
  sgdma_rx_csr_non_bursting_master_requests <= internal_cpuNios_data_master_requests_sgdma_rx_csr;
  --sgdma_rx_csr_any_bursting_master_saved_grant mux, which is an e_mux
  sgdma_rx_csr_any_bursting_master_saved_grant <= std_logic'('0');
  --sgdma_rx_csr_arb_share_counter_next_value assignment, which is an e_assign
  sgdma_rx_csr_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_rx_csr_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_rx_csr_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sgdma_rx_csr_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_rx_csr_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sgdma_rx_csr_allgrants all slave grants, which is an e_mux
  sgdma_rx_csr_allgrants <= sgdma_rx_csr_grant_vector;
  --sgdma_rx_csr_end_xfer assignment, which is an e_assign
  sgdma_rx_csr_end_xfer <= NOT ((sgdma_rx_csr_waits_for_read OR sgdma_rx_csr_waits_for_write));
  --end_xfer_arb_share_counter_term_sgdma_rx_csr arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sgdma_rx_csr <= sgdma_rx_csr_end_xfer AND (((NOT sgdma_rx_csr_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sgdma_rx_csr_arb_share_counter arbitration counter enable, which is an e_assign
  sgdma_rx_csr_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sgdma_rx_csr AND sgdma_rx_csr_allgrants)) OR ((end_xfer_arb_share_counter_term_sgdma_rx_csr AND NOT sgdma_rx_csr_non_bursting_master_requests));
  --sgdma_rx_csr_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_rx_csr_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sgdma_rx_csr_arb_counter_enable) = '1' then 
        sgdma_rx_csr_arb_share_counter <= sgdma_rx_csr_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sgdma_rx_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_rx_csr_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sgdma_rx_csr_master_qreq_vector AND end_xfer_arb_share_counter_term_sgdma_rx_csr)) OR ((end_xfer_arb_share_counter_term_sgdma_rx_csr AND NOT sgdma_rx_csr_non_bursting_master_requests)))) = '1' then 
        sgdma_rx_csr_slavearbiterlockenable <= sgdma_rx_csr_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master sgdma_rx/csr arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= sgdma_rx_csr_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --sgdma_rx_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sgdma_rx_csr_slavearbiterlockenable2 <= sgdma_rx_csr_arb_share_counter_next_value;
  --cpuNios/data_master sgdma_rx/csr arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= sgdma_rx_csr_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --sgdma_rx_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  sgdma_rx_csr_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_sgdma_rx_csr <= internal_cpuNios_data_master_requests_sgdma_rx_csr AND NOT (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write));
  --sgdma_rx_csr_writedata mux, which is an e_mux
  sgdma_rx_csr_writedata <= cpuNios_data_master_writedata;
  --master is always granted when requested
  internal_cpuNios_data_master_granted_sgdma_rx_csr <= internal_cpuNios_data_master_qualified_request_sgdma_rx_csr;
  --cpuNios/data_master saved-grant sgdma_rx/csr, which is an e_assign
  cpuNios_data_master_saved_grant_sgdma_rx_csr <= internal_cpuNios_data_master_requests_sgdma_rx_csr;
  --allow new arb cycle for sgdma_rx/csr, which is an e_assign
  sgdma_rx_csr_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sgdma_rx_csr_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sgdma_rx_csr_master_qreq_vector <= std_logic'('1');
  --sgdma_rx_csr_reset_n assignment, which is an e_assign
  sgdma_rx_csr_reset_n <= reset_n;
  sgdma_rx_csr_chipselect <= internal_cpuNios_data_master_granted_sgdma_rx_csr;
  --sgdma_rx_csr_firsttransfer first transaction, which is an e_assign
  sgdma_rx_csr_firsttransfer <= A_WE_StdLogic((std_logic'(sgdma_rx_csr_begins_xfer) = '1'), sgdma_rx_csr_unreg_firsttransfer, sgdma_rx_csr_reg_firsttransfer);
  --sgdma_rx_csr_unreg_firsttransfer first transaction, which is an e_assign
  sgdma_rx_csr_unreg_firsttransfer <= NOT ((sgdma_rx_csr_slavearbiterlockenable AND sgdma_rx_csr_any_continuerequest));
  --sgdma_rx_csr_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_rx_csr_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sgdma_rx_csr_begins_xfer) = '1' then 
        sgdma_rx_csr_reg_firsttransfer <= sgdma_rx_csr_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sgdma_rx_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sgdma_rx_csr_beginbursttransfer_internal <= sgdma_rx_csr_begins_xfer;
  --sgdma_rx_csr_read assignment, which is an e_mux
  sgdma_rx_csr_read <= internal_cpuNios_data_master_granted_sgdma_rx_csr AND cpuNios_data_master_read;
  --sgdma_rx_csr_write assignment, which is an e_mux
  sgdma_rx_csr_write <= internal_cpuNios_data_master_granted_sgdma_rx_csr AND cpuNios_data_master_write;
  shifted_address_to_sgdma_rx_csr_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --sgdma_rx_csr_address mux, which is an e_mux
  sgdma_rx_csr_address <= A_EXT (A_SRL(shifted_address_to_sgdma_rx_csr_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --d1_sgdma_rx_csr_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sgdma_rx_csr_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sgdma_rx_csr_end_xfer <= sgdma_rx_csr_end_xfer;
    end if;

  end process;

  --sgdma_rx_csr_waits_for_read in a cycle, which is an e_mux
  sgdma_rx_csr_waits_for_read <= sgdma_rx_csr_in_a_read_cycle AND sgdma_rx_csr_begins_xfer;
  --sgdma_rx_csr_in_a_read_cycle assignment, which is an e_assign
  sgdma_rx_csr_in_a_read_cycle <= internal_cpuNios_data_master_granted_sgdma_rx_csr AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sgdma_rx_csr_in_a_read_cycle;
  --sgdma_rx_csr_waits_for_write in a cycle, which is an e_mux
  sgdma_rx_csr_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_rx_csr_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sgdma_rx_csr_in_a_write_cycle assignment, which is an e_assign
  sgdma_rx_csr_in_a_write_cycle <= internal_cpuNios_data_master_granted_sgdma_rx_csr AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sgdma_rx_csr_in_a_write_cycle;
  wait_for_sgdma_rx_csr_counter <= std_logic'('0');
  --assign sgdma_rx_csr_irq_from_sa = sgdma_rx_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sgdma_rx_csr_irq_from_sa <= sgdma_rx_csr_irq;
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_sgdma_rx_csr <= internal_cpuNios_data_master_granted_sgdma_rx_csr;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_sgdma_rx_csr <= internal_cpuNios_data_master_qualified_request_sgdma_rx_csr;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_sgdma_rx_csr <= internal_cpuNios_data_master_requests_sgdma_rx_csr;
--synthesis translate_off
    --sgdma_rx/csr enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sgdma_rx_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_in_ready : IN STD_LOGIC;
                 signal tse_mac_receive_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_receive_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal tse_mac_receive_endofpacket : IN STD_LOGIC;
                 signal tse_mac_receive_error : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal tse_mac_receive_startofpacket : IN STD_LOGIC;
                 signal tse_mac_receive_valid : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_rx_in_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_in_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sgdma_rx_in_endofpacket : OUT STD_LOGIC;
                 signal sgdma_rx_in_error : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal sgdma_rx_in_ready_from_sa : OUT STD_LOGIC;
                 signal sgdma_rx_in_startofpacket : OUT STD_LOGIC;
                 signal sgdma_rx_in_valid : OUT STD_LOGIC
              );
end entity sgdma_rx_in_arbitrator;


architecture europa of sgdma_rx_in_arbitrator is

begin

  --mux sgdma_rx_in_data, which is an e_mux
  sgdma_rx_in_data <= tse_mac_receive_data;
  --mux sgdma_rx_in_empty, which is an e_mux
  sgdma_rx_in_empty <= tse_mac_receive_empty;
  --mux sgdma_rx_in_endofpacket, which is an e_mux
  sgdma_rx_in_endofpacket <= tse_mac_receive_endofpacket;
  --mux sgdma_rx_in_error, which is an e_mux
  sgdma_rx_in_error <= tse_mac_receive_error;
  --assign sgdma_rx_in_ready_from_sa = sgdma_rx_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  sgdma_rx_in_ready_from_sa <= sgdma_rx_in_ready;
  --mux sgdma_rx_in_startofpacket, which is an e_mux
  sgdma_rx_in_startofpacket <= tse_mac_receive_startofpacket;
  --mux sgdma_rx_in_valid, which is an e_mux
  sgdma_rx_in_valid <= tse_mac_receive_valid;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module;


architecture europa of selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_rx_descriptor_read_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_descriptor_offset_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal descriptor_offset_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (255 DOWNTO 0);
                 signal descriptor_offset_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_read : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_rx_descriptor_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_read_latency_counter : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_read_readdatavalid : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_rx_descriptor_read_arbitrator;


architecture europa of sgdma_rx_descriptor_read_arbitrator is
component selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module;

                signal active_and_waiting_last_time :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_readdata_from_sa_part_selected_by_negative_dbs :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal empty_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo :  STD_LOGIC;
                signal full_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_rx_descriptor_read_latency_counter :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_read_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal module_input31 :  STD_LOGIC;
                signal module_input32 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal module_input33 :  STD_LOGIC;
                signal p1_sgdma_rx_descriptor_read_latency_counter :  STD_LOGIC;
                signal pre_flush_sgdma_rx_descriptor_read_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal read_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo :  STD_LOGIC;
                signal selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sgdma_rx_descriptor_read_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_read_is_granted_some_slave :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read_but_no_slave_selected :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read_last_time :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_run :  STD_LOGIC;
                signal write_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 OR NOT sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 OR NOT sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 OR NOT (sgdma_rx_descriptor_read_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT descriptor_offset_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_rx_descriptor_read_read))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_rx_descriptor_read_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_rx_descriptor_read_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("00000") & sgdma_rx_descriptor_read_address(26 DOWNTO 0));
  --sgdma_rx_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_rx_descriptor_read_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      sgdma_rx_descriptor_read_read_but_no_slave_selected <= (sgdma_rx_descriptor_read_read AND sgdma_rx_descriptor_read_run) AND NOT sgdma_rx_descriptor_read_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  sgdma_rx_descriptor_read_is_granted_some_slave <= sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_sgdma_rx_descriptor_read_readdatavalid <= sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  sgdma_rx_descriptor_read_readdatavalid <= sgdma_rx_descriptor_read_read_but_no_slave_selected OR pre_flush_sgdma_rx_descriptor_read_readdatavalid;
  --Negative Dynamic Bus-sizing mux.
  --this mux selects the correct eighth of the 
  --wide data coming from the slave descriptor_offset_bridge/s1 
  descriptor_offset_bridge_s1_readdata_from_sa_part_selected_by_negative_dbs <= A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000000"))), descriptor_offset_bridge_s1_readdata_from_sa(31 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000001"))), descriptor_offset_bridge_s1_readdata_from_sa(63 DOWNTO 32), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000010"))), descriptor_offset_bridge_s1_readdata_from_sa(95 DOWNTO 64), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000011"))), descriptor_offset_bridge_s1_readdata_from_sa(127 DOWNTO 96), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000100"))), descriptor_offset_bridge_s1_readdata_from_sa(159 DOWNTO 128), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000101"))), descriptor_offset_bridge_s1_readdata_from_sa(191 DOWNTO 160), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000110"))), descriptor_offset_bridge_s1_readdata_from_sa(223 DOWNTO 192), descriptor_offset_bridge_s1_readdata_from_sa(255 DOWNTO 224))))))));
  --read_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo fifo read, which is an e_mux
  read_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo <= sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1;
  --write_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo fifo write, which is an e_mux
  write_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo <= (sgdma_rx_descriptor_read_read AND sgdma_rx_descriptor_read_run) AND sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1;
  selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1 <= selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output;
  --selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo, which is an e_fifo_with_registered_outputs
  selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo : selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module
    port map(
      data_out => selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output,
      empty => empty_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo,
      fifo_contains_ones_n => open,
      full => full_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo,
      clear_fifo => module_input31,
      clk => clk,
      data_in => module_input32,
      read => read_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo,
      reset_n => reset_n,
      sync_reset => module_input33,
      write => write_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo
    );

  module_input31 <= std_logic'('0');
  module_input32 <= internal_sgdma_rx_descriptor_read_address_to_slave(4 DOWNTO 2);
  module_input33 <= std_logic'('0');

  --sgdma_rx/descriptor_read readdata mux, which is an e_mux
  sgdma_rx_descriptor_read_readdata <= descriptor_offset_bridge_s1_readdata_from_sa_part_selected_by_negative_dbs;
  --actual waitrequest port, which is an e_assign
  internal_sgdma_rx_descriptor_read_waitrequest <= NOT sgdma_rx_descriptor_read_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_sgdma_rx_descriptor_read_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_sgdma_rx_descriptor_read_latency_counter <= p1_sgdma_rx_descriptor_read_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_sgdma_rx_descriptor_read_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((sgdma_rx_descriptor_read_run AND sgdma_rx_descriptor_read_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_read_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_sgdma_rx_descriptor_read_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_address_to_slave <= internal_sgdma_rx_descriptor_read_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_latency_counter <= internal_sgdma_rx_descriptor_read_latency_counter;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_waitrequest <= internal_sgdma_rx_descriptor_read_waitrequest;
--synthesis translate_off
    --sgdma_rx_descriptor_read_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_descriptor_read_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_rx_descriptor_read_address_last_time <= sgdma_rx_descriptor_read_address;
      end if;

    end process;

    --sgdma_rx/descriptor_read waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_rx_descriptor_read_waitrequest AND (sgdma_rx_descriptor_read_read);
      end if;

    end process;

    --sgdma_rx_descriptor_read_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line36 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_descriptor_read_address /= sgdma_rx_descriptor_read_address_last_time))))) = '1' then 
          write(write_line36, now);
          write(write_line36, string'(": "));
          write(write_line36, string'("sgdma_rx_descriptor_read_address did not heed wait!!!"));
          write(output, write_line36.all);
          deallocate (write_line36);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_descriptor_read_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_descriptor_read_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_rx_descriptor_read_read_last_time <= sgdma_rx_descriptor_read_read;
      end if;

    end process;

    --sgdma_rx_descriptor_read_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line37 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_rx_descriptor_read_read) /= std_logic'(sgdma_rx_descriptor_read_read_last_time)))))) = '1' then 
          write(write_line37, now);
          write(write_line37, string'(": "));
          write(write_line37, string'("sgdma_rx_descriptor_read_read did not heed wait!!!"));
          write(output, write_line37.all);
          deallocate (write_line37);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo read when empty, which is an e_process
    process (clk)
    VARIABLE write_line38 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((empty_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo AND read_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo)) = '1' then 
          write(write_line38, now);
          write(write_line38, string'(": "));
          write(write_line38, string'("sgdma_rx/descriptor_read negative rdv fifo selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo: read AND empty."));
          write(output, write_line38.all & CR);
          deallocate (write_line38);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo write when full, which is an e_process
    process (clk)
    VARIABLE write_line39 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((full_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo AND write_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo) AND NOT read_selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo)) = '1' then 
          write(write_line39, now);
          write(write_line39, string'(": "));
          write(write_line39, string'("sgdma_rx/descriptor_read negative rdv fifo selecto_nrdv_sgdma_rx_descriptor_read_3_descriptor_offset_bridge_s1_fifo: write AND full."));
          write(output, write_line39.all & CR);
          deallocate (write_line39);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_rx_descriptor_write_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_descriptor_offset_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal descriptor_offset_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_write : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal sgdma_rx_descriptor_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_write_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_rx_descriptor_write_arbitrator;


architecture europa of sgdma_rx_descriptor_write_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_rx_descriptor_write_waitrequest :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_write_run :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_write_last_time :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 OR NOT sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 OR NOT sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 OR NOT (sgdma_rx_descriptor_write_write))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT descriptor_offset_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_rx_descriptor_write_write))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_rx_descriptor_write_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_rx_descriptor_write_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("00000") & sgdma_rx_descriptor_write_address(26 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_sgdma_rx_descriptor_write_waitrequest <= NOT sgdma_rx_descriptor_write_run;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_write_address_to_slave <= internal_sgdma_rx_descriptor_write_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_write_waitrequest <= internal_sgdma_rx_descriptor_write_waitrequest;
--synthesis translate_off
    --sgdma_rx_descriptor_write_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_descriptor_write_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_rx_descriptor_write_address_last_time <= sgdma_rx_descriptor_write_address;
      end if;

    end process;

    --sgdma_rx/descriptor_write waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_rx_descriptor_write_waitrequest AND (sgdma_rx_descriptor_write_write);
      end if;

    end process;

    --sgdma_rx_descriptor_write_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line40 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_descriptor_write_address /= sgdma_rx_descriptor_write_address_last_time))))) = '1' then 
          write(write_line40, now);
          write(write_line40, string'(": "));
          write(write_line40, string'("sgdma_rx_descriptor_write_address did not heed wait!!!"));
          write(output, write_line40.all);
          deallocate (write_line40);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_descriptor_write_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_descriptor_write_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_rx_descriptor_write_write_last_time <= sgdma_rx_descriptor_write_write;
      end if;

    end process;

    --sgdma_rx_descriptor_write_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line41 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_rx_descriptor_write_write) /= std_logic'(sgdma_rx_descriptor_write_write_last_time)))))) = '1' then 
          write(write_line41, now);
          write(write_line41, string'(": "));
          write(write_line41, string'("sgdma_rx_descriptor_write_write did not heed wait!!!"));
          write(output, write_line41.all);
          deallocate (write_line41);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_descriptor_write_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_descriptor_write_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_rx_descriptor_write_writedata_last_time <= sgdma_rx_descriptor_write_writedata;
      end if;

    end process;

    --sgdma_rx_descriptor_write_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line42 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_descriptor_write_writedata /= sgdma_rx_descriptor_write_writedata_last_time)))) AND sgdma_rx_descriptor_write_write)) = '1' then 
          write(write_line42, now);
          write(write_line42, string'(": "));
          write(write_line42, string'("sgdma_rx_descriptor_write_writedata did not heed wait!!!"));
          write(output, write_line42.all);
          deallocate (write_line42);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_rx_m_write_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_tse_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_m_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_write : IN STD_LOGIC;
                 signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_rx_m_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_m_write_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_rx_m_write_arbitrator;


architecture europa of sgdma_rx_m_write_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_rx_m_write_waitrequest :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal sgdma_rx_m_write_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_m_write_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sgdma_rx_m_write_run :  STD_LOGIC;
                signal sgdma_rx_m_write_write_last_time :  STD_LOGIC;
                signal sgdma_rx_m_write_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 OR NOT sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 OR NOT sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 OR NOT (sgdma_rx_m_write_write))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT tse_ddr_clock_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_rx_m_write_write))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_rx_m_write_run <= r_2;
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_rx_m_write_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000000") & sgdma_rx_m_write_address(24 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_sgdma_rx_m_write_waitrequest <= NOT sgdma_rx_m_write_run;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_address_to_slave <= internal_sgdma_rx_m_write_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_waitrequest <= internal_sgdma_rx_m_write_waitrequest;
--synthesis translate_off
    --sgdma_rx_m_write_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_m_write_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_rx_m_write_address_last_time <= sgdma_rx_m_write_address;
      end if;

    end process;

    --sgdma_rx/m_write waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_rx_m_write_waitrequest AND (sgdma_rx_m_write_write);
      end if;

    end process;

    --sgdma_rx_m_write_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line43 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_m_write_address /= sgdma_rx_m_write_address_last_time))))) = '1' then 
          write(write_line43, now);
          write(write_line43, string'(": "));
          write(write_line43, string'("sgdma_rx_m_write_address did not heed wait!!!"));
          write(output, write_line43.all);
          deallocate (write_line43);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_m_write_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_m_write_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        sgdma_rx_m_write_byteenable_last_time <= sgdma_rx_m_write_byteenable;
      end if;

    end process;

    --sgdma_rx_m_write_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line44 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_m_write_byteenable /= sgdma_rx_m_write_byteenable_last_time))))) = '1' then 
          write(write_line44, now);
          write(write_line44, string'(": "));
          write(write_line44, string'("sgdma_rx_m_write_byteenable did not heed wait!!!"));
          write(output, write_line44.all);
          deallocate (write_line44);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_m_write_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_m_write_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_rx_m_write_write_last_time <= sgdma_rx_m_write_write;
      end if;

    end process;

    --sgdma_rx_m_write_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line45 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_rx_m_write_write) /= std_logic'(sgdma_rx_m_write_write_last_time)))))) = '1' then 
          write(write_line45, now);
          write(write_line45, string'(": "));
          write(write_line45, string'("sgdma_rx_m_write_write did not heed wait!!!"));
          write(output, write_line45.all);
          deallocate (write_line45);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_m_write_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_m_write_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_rx_m_write_writedata_last_time <= sgdma_rx_m_write_writedata;
      end if;

    end process;

    --sgdma_rx_m_write_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line46 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_m_write_writedata /= sgdma_rx_m_write_writedata_last_time)))) AND sgdma_rx_m_write_write)) = '1' then 
          write(write_line46, now);
          write(write_line46, string'(": "));
          write(write_line46, string'("sgdma_rx_m_write_writedata did not heed wait!!!"));
          write(output, write_line46.all);
          deallocate (write_line46);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sgdma_tx_csr_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_csr_irq : IN STD_LOGIC;
                 signal sgdma_tx_csr_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal cpuNios_data_master_granted_sgdma_tx_csr : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_sgdma_tx_csr : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_sgdma_tx_csr : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_sgdma_tx_csr : OUT STD_LOGIC;
                 signal d1_sgdma_tx_csr_end_xfer : OUT STD_LOGIC;
                 signal sgdma_tx_csr_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal sgdma_tx_csr_chipselect : OUT STD_LOGIC;
                 signal sgdma_tx_csr_irq_from_sa : OUT STD_LOGIC;
                 signal sgdma_tx_csr_read : OUT STD_LOGIC;
                 signal sgdma_tx_csr_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_csr_reset_n : OUT STD_LOGIC;
                 signal sgdma_tx_csr_write : OUT STD_LOGIC;
                 signal sgdma_tx_csr_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity sgdma_tx_csr_arbitrator;


architecture europa of sgdma_tx_csr_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_sgdma_tx_csr :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sgdma_tx_csr :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_sgdma_tx_csr :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_sgdma_tx_csr :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_sgdma_tx_csr :  STD_LOGIC;
                signal sgdma_tx_csr_allgrants :  STD_LOGIC;
                signal sgdma_tx_csr_allow_new_arb_cycle :  STD_LOGIC;
                signal sgdma_tx_csr_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sgdma_tx_csr_any_continuerequest :  STD_LOGIC;
                signal sgdma_tx_csr_arb_counter_enable :  STD_LOGIC;
                signal sgdma_tx_csr_arb_share_counter :  STD_LOGIC;
                signal sgdma_tx_csr_arb_share_counter_next_value :  STD_LOGIC;
                signal sgdma_tx_csr_arb_share_set_values :  STD_LOGIC;
                signal sgdma_tx_csr_beginbursttransfer_internal :  STD_LOGIC;
                signal sgdma_tx_csr_begins_xfer :  STD_LOGIC;
                signal sgdma_tx_csr_end_xfer :  STD_LOGIC;
                signal sgdma_tx_csr_firsttransfer :  STD_LOGIC;
                signal sgdma_tx_csr_grant_vector :  STD_LOGIC;
                signal sgdma_tx_csr_in_a_read_cycle :  STD_LOGIC;
                signal sgdma_tx_csr_in_a_write_cycle :  STD_LOGIC;
                signal sgdma_tx_csr_master_qreq_vector :  STD_LOGIC;
                signal sgdma_tx_csr_non_bursting_master_requests :  STD_LOGIC;
                signal sgdma_tx_csr_reg_firsttransfer :  STD_LOGIC;
                signal sgdma_tx_csr_slavearbiterlockenable :  STD_LOGIC;
                signal sgdma_tx_csr_slavearbiterlockenable2 :  STD_LOGIC;
                signal sgdma_tx_csr_unreg_firsttransfer :  STD_LOGIC;
                signal sgdma_tx_csr_waits_for_read :  STD_LOGIC;
                signal sgdma_tx_csr_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_sgdma_tx_csr_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal wait_for_sgdma_tx_csr_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sgdma_tx_csr_end_xfer;
    end if;

  end process;

  sgdma_tx_csr_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_sgdma_tx_csr);
  --assign sgdma_tx_csr_readdata_from_sa = sgdma_tx_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sgdma_tx_csr_readdata_from_sa <= sgdma_tx_csr_readdata;
  internal_cpuNios_data_master_requests_sgdma_tx_csr <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 6) & std_logic_vector'("000000")) = std_logic_vector'("100000000000100100101000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --sgdma_tx_csr_arb_share_counter set values, which is an e_mux
  sgdma_tx_csr_arb_share_set_values <= std_logic'('1');
  --sgdma_tx_csr_non_bursting_master_requests mux, which is an e_mux
  sgdma_tx_csr_non_bursting_master_requests <= internal_cpuNios_data_master_requests_sgdma_tx_csr;
  --sgdma_tx_csr_any_bursting_master_saved_grant mux, which is an e_mux
  sgdma_tx_csr_any_bursting_master_saved_grant <= std_logic'('0');
  --sgdma_tx_csr_arb_share_counter_next_value assignment, which is an e_assign
  sgdma_tx_csr_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_tx_csr_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_tx_csr_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sgdma_tx_csr_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_tx_csr_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sgdma_tx_csr_allgrants all slave grants, which is an e_mux
  sgdma_tx_csr_allgrants <= sgdma_tx_csr_grant_vector;
  --sgdma_tx_csr_end_xfer assignment, which is an e_assign
  sgdma_tx_csr_end_xfer <= NOT ((sgdma_tx_csr_waits_for_read OR sgdma_tx_csr_waits_for_write));
  --end_xfer_arb_share_counter_term_sgdma_tx_csr arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sgdma_tx_csr <= sgdma_tx_csr_end_xfer AND (((NOT sgdma_tx_csr_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sgdma_tx_csr_arb_share_counter arbitration counter enable, which is an e_assign
  sgdma_tx_csr_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sgdma_tx_csr AND sgdma_tx_csr_allgrants)) OR ((end_xfer_arb_share_counter_term_sgdma_tx_csr AND NOT sgdma_tx_csr_non_bursting_master_requests));
  --sgdma_tx_csr_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_csr_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sgdma_tx_csr_arb_counter_enable) = '1' then 
        sgdma_tx_csr_arb_share_counter <= sgdma_tx_csr_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sgdma_tx_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_csr_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sgdma_tx_csr_master_qreq_vector AND end_xfer_arb_share_counter_term_sgdma_tx_csr)) OR ((end_xfer_arb_share_counter_term_sgdma_tx_csr AND NOT sgdma_tx_csr_non_bursting_master_requests)))) = '1' then 
        sgdma_tx_csr_slavearbiterlockenable <= sgdma_tx_csr_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master sgdma_tx/csr arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= sgdma_tx_csr_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --sgdma_tx_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sgdma_tx_csr_slavearbiterlockenable2 <= sgdma_tx_csr_arb_share_counter_next_value;
  --cpuNios/data_master sgdma_tx/csr arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= sgdma_tx_csr_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --sgdma_tx_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  sgdma_tx_csr_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_sgdma_tx_csr <= internal_cpuNios_data_master_requests_sgdma_tx_csr AND NOT (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write));
  --sgdma_tx_csr_writedata mux, which is an e_mux
  sgdma_tx_csr_writedata <= cpuNios_data_master_writedata;
  --master is always granted when requested
  internal_cpuNios_data_master_granted_sgdma_tx_csr <= internal_cpuNios_data_master_qualified_request_sgdma_tx_csr;
  --cpuNios/data_master saved-grant sgdma_tx/csr, which is an e_assign
  cpuNios_data_master_saved_grant_sgdma_tx_csr <= internal_cpuNios_data_master_requests_sgdma_tx_csr;
  --allow new arb cycle for sgdma_tx/csr, which is an e_assign
  sgdma_tx_csr_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sgdma_tx_csr_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sgdma_tx_csr_master_qreq_vector <= std_logic'('1');
  --sgdma_tx_csr_reset_n assignment, which is an e_assign
  sgdma_tx_csr_reset_n <= reset_n;
  sgdma_tx_csr_chipselect <= internal_cpuNios_data_master_granted_sgdma_tx_csr;
  --sgdma_tx_csr_firsttransfer first transaction, which is an e_assign
  sgdma_tx_csr_firsttransfer <= A_WE_StdLogic((std_logic'(sgdma_tx_csr_begins_xfer) = '1'), sgdma_tx_csr_unreg_firsttransfer, sgdma_tx_csr_reg_firsttransfer);
  --sgdma_tx_csr_unreg_firsttransfer first transaction, which is an e_assign
  sgdma_tx_csr_unreg_firsttransfer <= NOT ((sgdma_tx_csr_slavearbiterlockenable AND sgdma_tx_csr_any_continuerequest));
  --sgdma_tx_csr_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_csr_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sgdma_tx_csr_begins_xfer) = '1' then 
        sgdma_tx_csr_reg_firsttransfer <= sgdma_tx_csr_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sgdma_tx_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sgdma_tx_csr_beginbursttransfer_internal <= sgdma_tx_csr_begins_xfer;
  --sgdma_tx_csr_read assignment, which is an e_mux
  sgdma_tx_csr_read <= internal_cpuNios_data_master_granted_sgdma_tx_csr AND cpuNios_data_master_read;
  --sgdma_tx_csr_write assignment, which is an e_mux
  sgdma_tx_csr_write <= internal_cpuNios_data_master_granted_sgdma_tx_csr AND cpuNios_data_master_write;
  shifted_address_to_sgdma_tx_csr_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --sgdma_tx_csr_address mux, which is an e_mux
  sgdma_tx_csr_address <= A_EXT (A_SRL(shifted_address_to_sgdma_tx_csr_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")), 4);
  --d1_sgdma_tx_csr_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sgdma_tx_csr_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sgdma_tx_csr_end_xfer <= sgdma_tx_csr_end_xfer;
    end if;

  end process;

  --sgdma_tx_csr_waits_for_read in a cycle, which is an e_mux
  sgdma_tx_csr_waits_for_read <= sgdma_tx_csr_in_a_read_cycle AND sgdma_tx_csr_begins_xfer;
  --sgdma_tx_csr_in_a_read_cycle assignment, which is an e_assign
  sgdma_tx_csr_in_a_read_cycle <= internal_cpuNios_data_master_granted_sgdma_tx_csr AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sgdma_tx_csr_in_a_read_cycle;
  --sgdma_tx_csr_waits_for_write in a cycle, which is an e_mux
  sgdma_tx_csr_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_tx_csr_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sgdma_tx_csr_in_a_write_cycle assignment, which is an e_assign
  sgdma_tx_csr_in_a_write_cycle <= internal_cpuNios_data_master_granted_sgdma_tx_csr AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sgdma_tx_csr_in_a_write_cycle;
  wait_for_sgdma_tx_csr_counter <= std_logic'('0');
  --assign sgdma_tx_csr_irq_from_sa = sgdma_tx_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sgdma_tx_csr_irq_from_sa <= sgdma_tx_csr_irq;
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_sgdma_tx_csr <= internal_cpuNios_data_master_granted_sgdma_tx_csr;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_sgdma_tx_csr <= internal_cpuNios_data_master_qualified_request_sgdma_tx_csr;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_sgdma_tx_csr <= internal_cpuNios_data_master_requests_sgdma_tx_csr;
--synthesis translate_off
    --sgdma_tx/csr enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module;


architecture europa of selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_0 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_1 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_2 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal stage_3 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_3;
  empty <= NOT(full_0);
  full_4 <= std_logic'('0');
  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic_vector'("000");
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic_vector'("000");
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic_vector'("000");
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic_vector'("000");
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(or_reduce(data_in)))), A_WE_StdLogicVector((std_logic'(((((read AND (or_reduce(data_in))) AND write) AND (or_reduce(stage_0))))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (or_reduce(data_in))))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (or_reduce(stage_0))))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_tx_descriptor_read_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_descriptor_offset_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal descriptor_offset_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (255 DOWNTO 0);
                 signal descriptor_offset_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_read : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_tx_descriptor_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_read_latency_counter : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_read_readdatavalid : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_tx_descriptor_read_arbitrator;


architecture europa of sgdma_tx_descriptor_read_arbitrator is
component selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module;

                signal active_and_waiting_last_time :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_readdata_from_sa_part_selected_by_negative_dbs :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal empty_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo :  STD_LOGIC;
                signal full_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_tx_descriptor_read_latency_counter :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_read_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal module_input34 :  STD_LOGIC;
                signal module_input35 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal module_input36 :  STD_LOGIC;
                signal p1_sgdma_tx_descriptor_read_latency_counter :  STD_LOGIC;
                signal pre_flush_sgdma_tx_descriptor_read_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal read_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo :  STD_LOGIC;
                signal selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1 :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sgdma_tx_descriptor_read_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_read_is_granted_some_slave :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read_but_no_slave_selected :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read_last_time :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_run :  STD_LOGIC;
                signal write_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 OR NOT sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 OR NOT sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 OR NOT (sgdma_tx_descriptor_read_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT descriptor_offset_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_tx_descriptor_read_read))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_tx_descriptor_read_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_tx_descriptor_read_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("00000") & sgdma_tx_descriptor_read_address(26 DOWNTO 0));
  --sgdma_tx_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_descriptor_read_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      sgdma_tx_descriptor_read_read_but_no_slave_selected <= (sgdma_tx_descriptor_read_read AND sgdma_tx_descriptor_read_run) AND NOT sgdma_tx_descriptor_read_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  sgdma_tx_descriptor_read_is_granted_some_slave <= sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_sgdma_tx_descriptor_read_readdatavalid <= sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  sgdma_tx_descriptor_read_readdatavalid <= sgdma_tx_descriptor_read_read_but_no_slave_selected OR pre_flush_sgdma_tx_descriptor_read_readdatavalid;
  --Negative Dynamic Bus-sizing mux.
  --this mux selects the correct eighth of the 
  --wide data coming from the slave descriptor_offset_bridge/s1 
  descriptor_offset_bridge_s1_readdata_from_sa_part_selected_by_negative_dbs <= A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000000"))), descriptor_offset_bridge_s1_readdata_from_sa(31 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000001"))), descriptor_offset_bridge_s1_readdata_from_sa(63 DOWNTO 32), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000010"))), descriptor_offset_bridge_s1_readdata_from_sa(95 DOWNTO 64), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000011"))), descriptor_offset_bridge_s1_readdata_from_sa(127 DOWNTO 96), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000100"))), descriptor_offset_bridge_s1_readdata_from_sa(159 DOWNTO 128), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000101"))), descriptor_offset_bridge_s1_readdata_from_sa(191 DOWNTO 160), A_WE_StdLogicVector((((std_logic_vector'("00000000000000000000000000000") & (selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1)) = std_logic_vector'("00000000000000000000000000000110"))), descriptor_offset_bridge_s1_readdata_from_sa(223 DOWNTO 192), descriptor_offset_bridge_s1_readdata_from_sa(255 DOWNTO 224))))))));
  --read_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo fifo read, which is an e_mux
  read_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo <= sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1;
  --write_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo fifo write, which is an e_mux
  write_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo <= (sgdma_tx_descriptor_read_read AND sgdma_tx_descriptor_read_run) AND sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1;
  selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output_descriptor_offset_bridge_s1 <= selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output;
  --selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo, which is an e_fifo_with_registered_outputs
  selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo : selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_module
    port map(
      data_out => selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo_output,
      empty => empty_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo,
      fifo_contains_ones_n => open,
      full => full_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo,
      clear_fifo => module_input34,
      clk => clk,
      data_in => module_input35,
      read => read_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo,
      reset_n => reset_n,
      sync_reset => module_input36,
      write => write_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo
    );

  module_input34 <= std_logic'('0');
  module_input35 <= internal_sgdma_tx_descriptor_read_address_to_slave(4 DOWNTO 2);
  module_input36 <= std_logic'('0');

  --sgdma_tx/descriptor_read readdata mux, which is an e_mux
  sgdma_tx_descriptor_read_readdata <= descriptor_offset_bridge_s1_readdata_from_sa_part_selected_by_negative_dbs;
  --actual waitrequest port, which is an e_assign
  internal_sgdma_tx_descriptor_read_waitrequest <= NOT sgdma_tx_descriptor_read_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_sgdma_tx_descriptor_read_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_sgdma_tx_descriptor_read_latency_counter <= p1_sgdma_tx_descriptor_read_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_sgdma_tx_descriptor_read_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((sgdma_tx_descriptor_read_run AND sgdma_tx_descriptor_read_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_sgdma_tx_descriptor_read_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_descriptor_read_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_address_to_slave <= internal_sgdma_tx_descriptor_read_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_latency_counter <= internal_sgdma_tx_descriptor_read_latency_counter;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_waitrequest <= internal_sgdma_tx_descriptor_read_waitrequest;
--synthesis translate_off
    --sgdma_tx_descriptor_read_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_descriptor_read_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_tx_descriptor_read_address_last_time <= sgdma_tx_descriptor_read_address;
      end if;

    end process;

    --sgdma_tx/descriptor_read waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_tx_descriptor_read_waitrequest AND (sgdma_tx_descriptor_read_read);
      end if;

    end process;

    --sgdma_tx_descriptor_read_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line47 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_tx_descriptor_read_address /= sgdma_tx_descriptor_read_address_last_time))))) = '1' then 
          write(write_line47, now);
          write(write_line47, string'(": "));
          write(write_line47, string'("sgdma_tx_descriptor_read_address did not heed wait!!!"));
          write(output, write_line47.all);
          deallocate (write_line47);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_tx_descriptor_read_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_descriptor_read_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_tx_descriptor_read_read_last_time <= sgdma_tx_descriptor_read_read;
      end if;

    end process;

    --sgdma_tx_descriptor_read_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line48 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_tx_descriptor_read_read) /= std_logic'(sgdma_tx_descriptor_read_read_last_time)))))) = '1' then 
          write(write_line48, now);
          write(write_line48, string'(": "));
          write(write_line48, string'("sgdma_tx_descriptor_read_read did not heed wait!!!"));
          write(output, write_line48.all);
          deallocate (write_line48);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo read when empty, which is an e_process
    process (clk)
    VARIABLE write_line49 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((empty_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo AND read_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo)) = '1' then 
          write(write_line49, now);
          write(write_line49, string'(": "));
          write(write_line49, string'("sgdma_tx/descriptor_read negative rdv fifo selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo: read AND empty."));
          write(output, write_line49.all & CR);
          deallocate (write_line49);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo write when full, which is an e_process
    process (clk)
    VARIABLE write_line50 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((full_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo AND write_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo) AND NOT read_selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo)) = '1' then 
          write(write_line50, now);
          write(write_line50, string'(": "));
          write(write_line50, string'("sgdma_tx/descriptor_read negative rdv fifo selecto_nrdv_sgdma_tx_descriptor_read_3_descriptor_offset_bridge_s1_fifo: write AND full."));
          write(output, write_line50.all & CR);
          deallocate (write_line50);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_tx_descriptor_write_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_descriptor_offset_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal descriptor_offset_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_write : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal sgdma_tx_descriptor_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_write_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_tx_descriptor_write_arbitrator;


architecture europa of sgdma_tx_descriptor_write_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_tx_descriptor_write_waitrequest :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_write_run :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_write_last_time :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 OR NOT sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 OR NOT sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 OR NOT (sgdma_tx_descriptor_write_write))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT descriptor_offset_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_tx_descriptor_write_write))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_tx_descriptor_write_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_tx_descriptor_write_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("00000") & sgdma_tx_descriptor_write_address(26 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_sgdma_tx_descriptor_write_waitrequest <= NOT sgdma_tx_descriptor_write_run;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_write_address_to_slave <= internal_sgdma_tx_descriptor_write_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_write_waitrequest <= internal_sgdma_tx_descriptor_write_waitrequest;
--synthesis translate_off
    --sgdma_tx_descriptor_write_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_descriptor_write_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_tx_descriptor_write_address_last_time <= sgdma_tx_descriptor_write_address;
      end if;

    end process;

    --sgdma_tx/descriptor_write waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_tx_descriptor_write_waitrequest AND (sgdma_tx_descriptor_write_write);
      end if;

    end process;

    --sgdma_tx_descriptor_write_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line51 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_tx_descriptor_write_address /= sgdma_tx_descriptor_write_address_last_time))))) = '1' then 
          write(write_line51, now);
          write(write_line51, string'(": "));
          write(write_line51, string'("sgdma_tx_descriptor_write_address did not heed wait!!!"));
          write(output, write_line51.all);
          deallocate (write_line51);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_tx_descriptor_write_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_descriptor_write_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_tx_descriptor_write_write_last_time <= sgdma_tx_descriptor_write_write;
      end if;

    end process;

    --sgdma_tx_descriptor_write_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line52 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_tx_descriptor_write_write) /= std_logic'(sgdma_tx_descriptor_write_write_last_time)))))) = '1' then 
          write(write_line52, now);
          write(write_line52, string'(": "));
          write(write_line52, string'("sgdma_tx_descriptor_write_write did not heed wait!!!"));
          write(output, write_line52.all);
          deallocate (write_line52);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_tx_descriptor_write_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_descriptor_write_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_tx_descriptor_write_writedata_last_time <= sgdma_tx_descriptor_write_writedata;
      end if;

    end process;

    --sgdma_tx_descriptor_write_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line53 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((sgdma_tx_descriptor_write_writedata /= sgdma_tx_descriptor_write_writedata_last_time)))) AND sgdma_tx_descriptor_write_write)) = '1' then 
          write(write_line53, now);
          write(write_line53, string'(": "));
          write(write_line53, string'("sgdma_tx_descriptor_write_writedata did not heed wait!!!"));
          write(output, write_line53.all);
          deallocate (write_line53);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_tx_m_read_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_tse_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_m_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1_shift_register : IN STD_LOGIC;
                 signal sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_tx_m_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_latency_counter : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_readdatavalid : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_tx_m_read_arbitrator;


architecture europa of sgdma_tx_m_read_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_tx_m_read_latency_counter :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_sgdma_tx_m_read_latency_counter :  STD_LOGIC;
                signal pre_flush_sgdma_tx_m_read_readdatavalid :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal sgdma_tx_m_read_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_m_read_is_granted_some_slave :  STD_LOGIC;
                signal sgdma_tx_m_read_read_but_no_slave_selected :  STD_LOGIC;
                signal sgdma_tx_m_read_read_last_time :  STD_LOGIC;
                signal sgdma_tx_m_read_run :  STD_LOGIC;

begin

  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 OR NOT sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 OR NOT sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 OR NOT (sgdma_tx_m_read_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT tse_ddr_clock_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_tx_m_read_read))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_tx_m_read_run <= r_2;
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_tx_m_read_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000000") & sgdma_tx_m_read_address(24 DOWNTO 0));
  --sgdma_tx_m_read_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_m_read_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      sgdma_tx_m_read_read_but_no_slave_selected <= (sgdma_tx_m_read_read AND sgdma_tx_m_read_run) AND NOT sgdma_tx_m_read_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  sgdma_tx_m_read_is_granted_some_slave <= sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_sgdma_tx_m_read_readdatavalid <= sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  sgdma_tx_m_read_readdatavalid <= sgdma_tx_m_read_read_but_no_slave_selected OR pre_flush_sgdma_tx_m_read_readdatavalid;
  --sgdma_tx/m_read readdata mux, which is an e_mux
  sgdma_tx_m_read_readdata <= tse_ddr_clock_bridge_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_sgdma_tx_m_read_waitrequest <= NOT sgdma_tx_m_read_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_sgdma_tx_m_read_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_sgdma_tx_m_read_latency_counter <= p1_sgdma_tx_m_read_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_sgdma_tx_m_read_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((sgdma_tx_m_read_run AND sgdma_tx_m_read_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_sgdma_tx_m_read_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_m_read_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --vhdl renameroo for output signals
  sgdma_tx_m_read_address_to_slave <= internal_sgdma_tx_m_read_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_latency_counter <= internal_sgdma_tx_m_read_latency_counter;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_waitrequest <= internal_sgdma_tx_m_read_waitrequest;
--synthesis translate_off
    --sgdma_tx_m_read_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_m_read_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_tx_m_read_address_last_time <= sgdma_tx_m_read_address;
      end if;

    end process;

    --sgdma_tx/m_read waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_tx_m_read_waitrequest AND (sgdma_tx_m_read_read);
      end if;

    end process;

    --sgdma_tx_m_read_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line54 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_tx_m_read_address /= sgdma_tx_m_read_address_last_time))))) = '1' then 
          write(write_line54, now);
          write(write_line54, string'(": "));
          write(write_line54, string'("sgdma_tx_m_read_address did not heed wait!!!"));
          write(output, write_line54.all);
          deallocate (write_line54);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_tx_m_read_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_m_read_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_tx_m_read_read_last_time <= sgdma_tx_m_read_read;
      end if;

    end process;

    --sgdma_tx_m_read_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line55 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_tx_m_read_read) /= std_logic'(sgdma_tx_m_read_read_last_time)))))) = '1' then 
          write(write_line55, now);
          write(write_line55, string'(": "));
          write(write_line55, string'("sgdma_tx_m_read_read did not heed wait!!!"));
          write(output, write_line55.all);
          deallocate (write_line55);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sgdma_tx_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sgdma_tx_out_endofpacket : IN STD_LOGIC;
                 signal sgdma_tx_out_error : IN STD_LOGIC;
                 signal sgdma_tx_out_startofpacket : IN STD_LOGIC;
                 signal sgdma_tx_out_valid : IN STD_LOGIC;
                 signal tse_mac_transmit_ready_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_tx_out_ready : OUT STD_LOGIC
              );
end entity sgdma_tx_out_arbitrator;


architecture europa of sgdma_tx_out_arbitrator is

begin

  --mux sgdma_tx_out_ready, which is an e_mux
  sgdma_tx_out_ready <= tse_mac_transmit_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sys_clk_timer_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_timer_s1_irq : IN STD_LOGIC;
                 signal sys_clk_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal cpuNios_data_master_granted_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal d1_sys_clk_timer_s1_end_xfer : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal sys_clk_timer_s1_chipselect : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_irq_from_sa : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sys_clk_timer_s1_reset_n : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_write_n : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sys_clk_timer_s1_arbitrator;


architecture europa of sys_clk_timer_s1_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_sys_clk_timer_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sys_clk_timer_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_sys_clk_timer_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_sys_clk_timer_s1 :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_sys_clk_timer_s1 :  STD_LOGIC;
                signal shifted_address_to_sys_clk_timer_s1_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal sys_clk_timer_s1_allgrants :  STD_LOGIC;
                signal sys_clk_timer_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sys_clk_timer_s1_any_continuerequest :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_counter_enable :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_share_counter :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_share_set_values :  STD_LOGIC;
                signal sys_clk_timer_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sys_clk_timer_s1_begins_xfer :  STD_LOGIC;
                signal sys_clk_timer_s1_end_xfer :  STD_LOGIC;
                signal sys_clk_timer_s1_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_grant_vector :  STD_LOGIC;
                signal sys_clk_timer_s1_in_a_read_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_in_a_write_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_master_qreq_vector :  STD_LOGIC;
                signal sys_clk_timer_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sys_clk_timer_s1_reg_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sys_clk_timer_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sys_clk_timer_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_waits_for_read :  STD_LOGIC;
                signal sys_clk_timer_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_sys_clk_timer_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sys_clk_timer_s1_end_xfer;
    end if;

  end process;

  sys_clk_timer_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_sys_clk_timer_s1);
  --assign sys_clk_timer_s1_readdata_from_sa = sys_clk_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sys_clk_timer_s1_readdata_from_sa <= sys_clk_timer_s1_readdata;
  internal_cpuNios_data_master_requests_sys_clk_timer_s1 <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("100000000000100011000000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --sys_clk_timer_s1_arb_share_counter set values, which is an e_mux
  sys_clk_timer_s1_arb_share_set_values <= std_logic'('1');
  --sys_clk_timer_s1_non_bursting_master_requests mux, which is an e_mux
  sys_clk_timer_s1_non_bursting_master_requests <= internal_cpuNios_data_master_requests_sys_clk_timer_s1;
  --sys_clk_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sys_clk_timer_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sys_clk_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  sys_clk_timer_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sys_clk_timer_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_timer_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sys_clk_timer_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_timer_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sys_clk_timer_s1_allgrants all slave grants, which is an e_mux
  sys_clk_timer_s1_allgrants <= sys_clk_timer_s1_grant_vector;
  --sys_clk_timer_s1_end_xfer assignment, which is an e_assign
  sys_clk_timer_s1_end_xfer <= NOT ((sys_clk_timer_s1_waits_for_read OR sys_clk_timer_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sys_clk_timer_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sys_clk_timer_s1 <= sys_clk_timer_s1_end_xfer AND (((NOT sys_clk_timer_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sys_clk_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sys_clk_timer_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND sys_clk_timer_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND NOT sys_clk_timer_s1_non_bursting_master_requests));
  --sys_clk_timer_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sys_clk_timer_s1_arb_counter_enable) = '1' then 
        sys_clk_timer_s1_arb_share_counter <= sys_clk_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sys_clk_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sys_clk_timer_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_sys_clk_timer_s1)) OR ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND NOT sys_clk_timer_s1_non_bursting_master_requests)))) = '1' then 
        sys_clk_timer_s1_slavearbiterlockenable <= sys_clk_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master sys_clk_timer/s1 arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= sys_clk_timer_s1_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --sys_clk_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sys_clk_timer_s1_slavearbiterlockenable2 <= sys_clk_timer_s1_arb_share_counter_next_value;
  --cpuNios/data_master sys_clk_timer/s1 arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= sys_clk_timer_s1_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --sys_clk_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  sys_clk_timer_s1_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_sys_clk_timer_s1 <= internal_cpuNios_data_master_requests_sys_clk_timer_s1 AND NOT (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write));
  --sys_clk_timer_s1_writedata mux, which is an e_mux
  sys_clk_timer_s1_writedata <= cpuNios_data_master_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_cpuNios_data_master_granted_sys_clk_timer_s1 <= internal_cpuNios_data_master_qualified_request_sys_clk_timer_s1;
  --cpuNios/data_master saved-grant sys_clk_timer/s1, which is an e_assign
  cpuNios_data_master_saved_grant_sys_clk_timer_s1 <= internal_cpuNios_data_master_requests_sys_clk_timer_s1;
  --allow new arb cycle for sys_clk_timer/s1, which is an e_assign
  sys_clk_timer_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sys_clk_timer_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sys_clk_timer_s1_master_qreq_vector <= std_logic'('1');
  --sys_clk_timer_s1_reset_n assignment, which is an e_assign
  sys_clk_timer_s1_reset_n <= reset_n;
  sys_clk_timer_s1_chipselect <= internal_cpuNios_data_master_granted_sys_clk_timer_s1;
  --sys_clk_timer_s1_firsttransfer first transaction, which is an e_assign
  sys_clk_timer_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sys_clk_timer_s1_begins_xfer) = '1'), sys_clk_timer_s1_unreg_firsttransfer, sys_clk_timer_s1_reg_firsttransfer);
  --sys_clk_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  sys_clk_timer_s1_unreg_firsttransfer <= NOT ((sys_clk_timer_s1_slavearbiterlockenable AND sys_clk_timer_s1_any_continuerequest));
  --sys_clk_timer_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sys_clk_timer_s1_begins_xfer) = '1' then 
        sys_clk_timer_s1_reg_firsttransfer <= sys_clk_timer_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sys_clk_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sys_clk_timer_s1_beginbursttransfer_internal <= sys_clk_timer_s1_begins_xfer;
  --~sys_clk_timer_s1_write_n assignment, which is an e_mux
  sys_clk_timer_s1_write_n <= NOT ((internal_cpuNios_data_master_granted_sys_clk_timer_s1 AND cpuNios_data_master_write));
  shifted_address_to_sys_clk_timer_s1_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --sys_clk_timer_s1_address mux, which is an e_mux
  sys_clk_timer_s1_address <= A_EXT (A_SRL(shifted_address_to_sys_clk_timer_s1_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_sys_clk_timer_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sys_clk_timer_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sys_clk_timer_s1_end_xfer <= sys_clk_timer_s1_end_xfer;
    end if;

  end process;

  --sys_clk_timer_s1_waits_for_read in a cycle, which is an e_mux
  sys_clk_timer_s1_waits_for_read <= sys_clk_timer_s1_in_a_read_cycle AND sys_clk_timer_s1_begins_xfer;
  --sys_clk_timer_s1_in_a_read_cycle assignment, which is an e_assign
  sys_clk_timer_s1_in_a_read_cycle <= internal_cpuNios_data_master_granted_sys_clk_timer_s1 AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sys_clk_timer_s1_in_a_read_cycle;
  --sys_clk_timer_s1_waits_for_write in a cycle, which is an e_mux
  sys_clk_timer_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_timer_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sys_clk_timer_s1_in_a_write_cycle assignment, which is an e_assign
  sys_clk_timer_s1_in_a_write_cycle <= internal_cpuNios_data_master_granted_sys_clk_timer_s1 AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sys_clk_timer_s1_in_a_write_cycle;
  wait_for_sys_clk_timer_s1_counter <= std_logic'('0');
  --assign sys_clk_timer_s1_irq_from_sa = sys_clk_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sys_clk_timer_s1_irq_from_sa <= sys_clk_timer_s1_irq;
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_sys_clk_timer_s1 <= internal_cpuNios_data_master_granted_sys_clk_timer_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_sys_clk_timer_s1 <= internal_cpuNios_data_master_qualified_request_sys_clk_timer_s1;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_sys_clk_timer_s1 <= internal_cpuNios_data_master_requests_sys_clk_timer_s1;
--synthesis translate_off
    --sys_clk_timer/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sysid_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal cpuNios_data_master_granted_sysid_control_slave : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_sysid_control_slave : OUT STD_LOGIC;
                 signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                 signal sysid_control_slave_address : OUT STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sysid_control_slave_reset_n : OUT STD_LOGIC
              );
end entity sysid_control_slave_arbitrator;


architecture europa of sysid_control_slave_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_sysid_control_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sysid_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_sysid_control_slave :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_sysid_control_slave :  STD_LOGIC;
                signal shifted_address_to_sysid_control_slave_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal sysid_control_slave_allgrants :  STD_LOGIC;
                signal sysid_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal sysid_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sysid_control_slave_any_continuerequest :  STD_LOGIC;
                signal sysid_control_slave_arb_counter_enable :  STD_LOGIC;
                signal sysid_control_slave_arb_share_counter :  STD_LOGIC;
                signal sysid_control_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal sysid_control_slave_arb_share_set_values :  STD_LOGIC;
                signal sysid_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal sysid_control_slave_begins_xfer :  STD_LOGIC;
                signal sysid_control_slave_end_xfer :  STD_LOGIC;
                signal sysid_control_slave_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_grant_vector :  STD_LOGIC;
                signal sysid_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal sysid_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal sysid_control_slave_master_qreq_vector :  STD_LOGIC;
                signal sysid_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal sysid_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal sysid_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_waits_for_read :  STD_LOGIC;
                signal sysid_control_slave_waits_for_write :  STD_LOGIC;
                signal wait_for_sysid_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sysid_control_slave_end_xfer;
    end if;

  end process;

  sysid_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_sysid_control_slave);
  --assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sysid_control_slave_readdata_from_sa <= sysid_control_slave_readdata;
  internal_cpuNios_data_master_requests_sysid_control_slave <= ((to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("100000000000100100011000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write)))) AND cpuNios_data_master_read;
  --sysid_control_slave_arb_share_counter set values, which is an e_mux
  sysid_control_slave_arb_share_set_values <= std_logic'('1');
  --sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  sysid_control_slave_non_bursting_master_requests <= internal_cpuNios_data_master_requests_sysid_control_slave;
  --sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  sysid_control_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  sysid_control_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sysid_control_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sysid_control_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sysid_control_slave_allgrants all slave grants, which is an e_mux
  sysid_control_slave_allgrants <= sysid_control_slave_grant_vector;
  --sysid_control_slave_end_xfer assignment, which is an e_assign
  sysid_control_slave_end_xfer <= NOT ((sysid_control_slave_waits_for_read OR sysid_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sysid_control_slave <= sysid_control_slave_end_xfer AND (((NOT sysid_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  sysid_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sysid_control_slave AND sysid_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests));
  --sysid_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_arb_counter_enable) = '1' then 
        sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sysid_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_sysid_control_slave)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests)))) = '1' then 
        sysid_control_slave_slavearbiterlockenable <= sysid_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master sysid/control_slave arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= sysid_control_slave_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sysid_control_slave_slavearbiterlockenable2 <= sysid_control_slave_arb_share_counter_next_value;
  --cpuNios/data_master sysid/control_slave arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= sysid_control_slave_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  sysid_control_slave_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_sysid_control_slave <= internal_cpuNios_data_master_requests_sysid_control_slave;
  --master is always granted when requested
  internal_cpuNios_data_master_granted_sysid_control_slave <= internal_cpuNios_data_master_qualified_request_sysid_control_slave;
  --cpuNios/data_master saved-grant sysid/control_slave, which is an e_assign
  cpuNios_data_master_saved_grant_sysid_control_slave <= internal_cpuNios_data_master_requests_sysid_control_slave;
  --allow new arb cycle for sysid/control_slave, which is an e_assign
  sysid_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sysid_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sysid_control_slave_master_qreq_vector <= std_logic'('1');
  --sysid_control_slave_reset_n assignment, which is an e_assign
  sysid_control_slave_reset_n <= reset_n;
  --sysid_control_slave_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(sysid_control_slave_begins_xfer) = '1'), sysid_control_slave_unreg_firsttransfer, sysid_control_slave_reg_firsttransfer);
  --sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_unreg_firsttransfer <= NOT ((sysid_control_slave_slavearbiterlockenable AND sysid_control_slave_any_continuerequest));
  --sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_begins_xfer) = '1' then 
        sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sysid_control_slave_beginbursttransfer_internal <= sysid_control_slave_begins_xfer;
  shifted_address_to_sysid_control_slave_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --sysid_control_slave_address mux, which is an e_mux
  sysid_control_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_sysid_control_slave_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_sysid_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sysid_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end if;

  end process;

  --sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  sysid_control_slave_waits_for_read <= sysid_control_slave_in_a_read_cycle AND sysid_control_slave_begins_xfer;
  --sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_read_cycle <= internal_cpuNios_data_master_granted_sysid_control_slave AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sysid_control_slave_in_a_read_cycle;
  --sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  sysid_control_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_write_cycle <= internal_cpuNios_data_master_granted_sysid_control_slave AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sysid_control_slave_in_a_write_cycle;
  wait_for_sysid_control_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_sysid_control_slave <= internal_cpuNios_data_master_granted_sysid_control_slave;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_sysid_control_slave <= internal_cpuNios_data_master_qualified_request_sysid_control_slave;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_sysid_control_slave <= internal_cpuNios_data_master_requests_sysid_control_slave;
--synthesis translate_off
    --sysid/control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_sgdma_tx_m_read_to_tse_ddr_clock_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_sgdma_tx_m_read_to_tse_ddr_clock_bridge_s1_module;


architecture europa of rdv_fifo_for_sgdma_tx_m_read_to_tse_ddr_clock_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_33 :  STD_LOGIC;
                signal full_34 :  STD_LOGIC;
                signal full_35 :  STD_LOGIC;
                signal full_36 :  STD_LOGIC;
                signal full_37 :  STD_LOGIC;
                signal full_38 :  STD_LOGIC;
                signal full_39 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_40 :  STD_LOGIC;
                signal full_41 :  STD_LOGIC;
                signal full_42 :  STD_LOGIC;
                signal full_43 :  STD_LOGIC;
                signal full_44 :  STD_LOGIC;
                signal full_45 :  STD_LOGIC;
                signal full_46 :  STD_LOGIC;
                signal full_47 :  STD_LOGIC;
                signal full_48 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p32_full_32 :  STD_LOGIC;
                signal p32_stage_32 :  STD_LOGIC;
                signal p33_full_33 :  STD_LOGIC;
                signal p33_stage_33 :  STD_LOGIC;
                signal p34_full_34 :  STD_LOGIC;
                signal p34_stage_34 :  STD_LOGIC;
                signal p35_full_35 :  STD_LOGIC;
                signal p35_stage_35 :  STD_LOGIC;
                signal p36_full_36 :  STD_LOGIC;
                signal p36_stage_36 :  STD_LOGIC;
                signal p37_full_37 :  STD_LOGIC;
                signal p37_stage_37 :  STD_LOGIC;
                signal p38_full_38 :  STD_LOGIC;
                signal p38_stage_38 :  STD_LOGIC;
                signal p39_full_39 :  STD_LOGIC;
                signal p39_stage_39 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p40_full_40 :  STD_LOGIC;
                signal p40_stage_40 :  STD_LOGIC;
                signal p41_full_41 :  STD_LOGIC;
                signal p41_stage_41 :  STD_LOGIC;
                signal p42_full_42 :  STD_LOGIC;
                signal p42_stage_42 :  STD_LOGIC;
                signal p43_full_43 :  STD_LOGIC;
                signal p43_stage_43 :  STD_LOGIC;
                signal p44_full_44 :  STD_LOGIC;
                signal p44_stage_44 :  STD_LOGIC;
                signal p45_full_45 :  STD_LOGIC;
                signal p45_stage_45 :  STD_LOGIC;
                signal p46_full_46 :  STD_LOGIC;
                signal p46_stage_46 :  STD_LOGIC;
                signal p47_full_47 :  STD_LOGIC;
                signal p47_stage_47 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_32 :  STD_LOGIC;
                signal stage_33 :  STD_LOGIC;
                signal stage_34 :  STD_LOGIC;
                signal stage_35 :  STD_LOGIC;
                signal stage_36 :  STD_LOGIC;
                signal stage_37 :  STD_LOGIC;
                signal stage_38 :  STD_LOGIC;
                signal stage_39 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_40 :  STD_LOGIC;
                signal stage_41 :  STD_LOGIC;
                signal stage_42 :  STD_LOGIC;
                signal stage_43 :  STD_LOGIC;
                signal stage_44 :  STD_LOGIC;
                signal stage_45 :  STD_LOGIC;
                signal stage_46 :  STD_LOGIC;
                signal stage_47 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_47;
  empty <= NOT(full_0);
  full_48 <= std_logic'('0');
  --data_47, which is an e_mux
  p47_stage_47 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_48 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_47, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_47 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_47))))) = '1' then 
        if std_logic'(((sync_reset AND full_47) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_48))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_47 <= std_logic'('0');
        else
          stage_47 <= p47_stage_47;
        end if;
      end if;
    end if;

  end process;

  --control_47, which is an e_mux
  p47_full_47 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_46))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_47, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_47 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_47 <= std_logic'('0');
        else
          full_47 <= p47_full_47;
        end if;
      end if;
    end if;

  end process;

  --data_46, which is an e_mux
  p46_stage_46 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_47 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_47);
  --data_reg_46, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_46 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_46))))) = '1' then 
        if std_logic'(((sync_reset AND full_46) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_47))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_46 <= std_logic'('0');
        else
          stage_46 <= p46_stage_46;
        end if;
      end if;
    end if;

  end process;

  --control_46, which is an e_mux
  p46_full_46 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_45, full_47);
  --control_reg_46, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_46 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_46 <= std_logic'('0');
        else
          full_46 <= p46_full_46;
        end if;
      end if;
    end if;

  end process;

  --data_45, which is an e_mux
  p45_stage_45 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_46 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_46);
  --data_reg_45, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_45 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_45))))) = '1' then 
        if std_logic'(((sync_reset AND full_45) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_46))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_45 <= std_logic'('0');
        else
          stage_45 <= p45_stage_45;
        end if;
      end if;
    end if;

  end process;

  --control_45, which is an e_mux
  p45_full_45 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_44, full_46);
  --control_reg_45, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_45 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_45 <= std_logic'('0');
        else
          full_45 <= p45_full_45;
        end if;
      end if;
    end if;

  end process;

  --data_44, which is an e_mux
  p44_stage_44 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_45 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_45);
  --data_reg_44, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_44 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_44))))) = '1' then 
        if std_logic'(((sync_reset AND full_44) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_45))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_44 <= std_logic'('0');
        else
          stage_44 <= p44_stage_44;
        end if;
      end if;
    end if;

  end process;

  --control_44, which is an e_mux
  p44_full_44 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_43, full_45);
  --control_reg_44, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_44 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_44 <= std_logic'('0');
        else
          full_44 <= p44_full_44;
        end if;
      end if;
    end if;

  end process;

  --data_43, which is an e_mux
  p43_stage_43 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_44 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_44);
  --data_reg_43, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_43 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_43))))) = '1' then 
        if std_logic'(((sync_reset AND full_43) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_44))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_43 <= std_logic'('0');
        else
          stage_43 <= p43_stage_43;
        end if;
      end if;
    end if;

  end process;

  --control_43, which is an e_mux
  p43_full_43 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_42, full_44);
  --control_reg_43, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_43 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_43 <= std_logic'('0');
        else
          full_43 <= p43_full_43;
        end if;
      end if;
    end if;

  end process;

  --data_42, which is an e_mux
  p42_stage_42 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_43 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_43);
  --data_reg_42, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_42 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_42))))) = '1' then 
        if std_logic'(((sync_reset AND full_42) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_43))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_42 <= std_logic'('0');
        else
          stage_42 <= p42_stage_42;
        end if;
      end if;
    end if;

  end process;

  --control_42, which is an e_mux
  p42_full_42 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_41, full_43);
  --control_reg_42, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_42 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_42 <= std_logic'('0');
        else
          full_42 <= p42_full_42;
        end if;
      end if;
    end if;

  end process;

  --data_41, which is an e_mux
  p41_stage_41 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_42 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_42);
  --data_reg_41, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_41 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_41))))) = '1' then 
        if std_logic'(((sync_reset AND full_41) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_42))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_41 <= std_logic'('0');
        else
          stage_41 <= p41_stage_41;
        end if;
      end if;
    end if;

  end process;

  --control_41, which is an e_mux
  p41_full_41 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_40, full_42);
  --control_reg_41, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_41 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_41 <= std_logic'('0');
        else
          full_41 <= p41_full_41;
        end if;
      end if;
    end if;

  end process;

  --data_40, which is an e_mux
  p40_stage_40 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_41 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_41);
  --data_reg_40, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_40 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_40))))) = '1' then 
        if std_logic'(((sync_reset AND full_40) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_41))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_40 <= std_logic'('0');
        else
          stage_40 <= p40_stage_40;
        end if;
      end if;
    end if;

  end process;

  --control_40, which is an e_mux
  p40_full_40 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_39, full_41);
  --control_reg_40, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_40 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_40 <= std_logic'('0');
        else
          full_40 <= p40_full_40;
        end if;
      end if;
    end if;

  end process;

  --data_39, which is an e_mux
  p39_stage_39 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_40 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_40);
  --data_reg_39, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_39 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_39))))) = '1' then 
        if std_logic'(((sync_reset AND full_39) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_40))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_39 <= std_logic'('0');
        else
          stage_39 <= p39_stage_39;
        end if;
      end if;
    end if;

  end process;

  --control_39, which is an e_mux
  p39_full_39 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_38, full_40);
  --control_reg_39, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_39 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_39 <= std_logic'('0');
        else
          full_39 <= p39_full_39;
        end if;
      end if;
    end if;

  end process;

  --data_38, which is an e_mux
  p38_stage_38 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_39 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_39);
  --data_reg_38, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_38 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_38))))) = '1' then 
        if std_logic'(((sync_reset AND full_38) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_39))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_38 <= std_logic'('0');
        else
          stage_38 <= p38_stage_38;
        end if;
      end if;
    end if;

  end process;

  --control_38, which is an e_mux
  p38_full_38 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_37, full_39);
  --control_reg_38, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_38 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_38 <= std_logic'('0');
        else
          full_38 <= p38_full_38;
        end if;
      end if;
    end if;

  end process;

  --data_37, which is an e_mux
  p37_stage_37 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_38 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_38);
  --data_reg_37, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_37 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_37))))) = '1' then 
        if std_logic'(((sync_reset AND full_37) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_38))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_37 <= std_logic'('0');
        else
          stage_37 <= p37_stage_37;
        end if;
      end if;
    end if;

  end process;

  --control_37, which is an e_mux
  p37_full_37 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_36, full_38);
  --control_reg_37, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_37 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_37 <= std_logic'('0');
        else
          full_37 <= p37_full_37;
        end if;
      end if;
    end if;

  end process;

  --data_36, which is an e_mux
  p36_stage_36 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_37 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_37);
  --data_reg_36, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_36 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_36))))) = '1' then 
        if std_logic'(((sync_reset AND full_36) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_37))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_36 <= std_logic'('0');
        else
          stage_36 <= p36_stage_36;
        end if;
      end if;
    end if;

  end process;

  --control_36, which is an e_mux
  p36_full_36 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_35, full_37);
  --control_reg_36, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_36 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_36 <= std_logic'('0');
        else
          full_36 <= p36_full_36;
        end if;
      end if;
    end if;

  end process;

  --data_35, which is an e_mux
  p35_stage_35 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_36 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_36);
  --data_reg_35, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_35 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_35))))) = '1' then 
        if std_logic'(((sync_reset AND full_35) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_36))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_35 <= std_logic'('0');
        else
          stage_35 <= p35_stage_35;
        end if;
      end if;
    end if;

  end process;

  --control_35, which is an e_mux
  p35_full_35 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_34, full_36);
  --control_reg_35, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_35 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_35 <= std_logic'('0');
        else
          full_35 <= p35_full_35;
        end if;
      end if;
    end if;

  end process;

  --data_34, which is an e_mux
  p34_stage_34 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_35 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_35);
  --data_reg_34, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_34 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_34))))) = '1' then 
        if std_logic'(((sync_reset AND full_34) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_35))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_34 <= std_logic'('0');
        else
          stage_34 <= p34_stage_34;
        end if;
      end if;
    end if;

  end process;

  --control_34, which is an e_mux
  p34_full_34 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_33, full_35);
  --control_reg_34, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_34 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_34 <= std_logic'('0');
        else
          full_34 <= p34_full_34;
        end if;
      end if;
    end if;

  end process;

  --data_33, which is an e_mux
  p33_stage_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_34 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_34);
  --data_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_33))))) = '1' then 
        if std_logic'(((sync_reset AND full_33) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_34))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_33 <= std_logic'('0');
        else
          stage_33 <= p33_stage_33;
        end if;
      end if;
    end if;

  end process;

  --control_33, which is an e_mux
  p33_full_33 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_32, full_34);
  --control_reg_33, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_33 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_33 <= std_logic'('0');
        else
          full_33 <= p33_full_33;
        end if;
      end if;
    end if;

  end process;

  --data_32, which is an e_mux
  p32_stage_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_33 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_33);
  --data_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_32))))) = '1' then 
        if std_logic'(((sync_reset AND full_32) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_33))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_32 <= std_logic'('0');
        else
          stage_32 <= p32_stage_32;
        end if;
      end if;
    end if;

  end process;

  --control_32, which is an e_mux
  p32_full_32 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_31, full_33);
  --control_reg_32, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_32 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_32 <= std_logic'('0');
        else
          full_32 <= p32_full_32;
        end if;
      end if;
    end if;

  end process;

  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_32);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_30, full_32);
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity tse_ddr_clock_bridge_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_m_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal sgdma_rx_m_write_write : IN STD_LOGIC;
                 signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_latency_counter : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_s1_endofpacket : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_ddr_clock_bridge_s1_readdatavalid : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_s1_waitrequest : IN STD_LOGIC;

              -- outputs:
                 signal d1_tse_ddr_clock_bridge_s1_end_xfer : OUT STD_LOGIC;
                 signal sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal tse_ddr_clock_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal tse_ddr_clock_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal tse_ddr_clock_bridge_s1_read : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_ddr_clock_bridge_s1_reset_n : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_s1_write : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity tse_ddr_clock_bridge_s1_arbitrator;


architecture europa of tse_ddr_clock_bridge_s1_arbitrator is
component rdv_fifo_for_sgdma_tx_m_read_to_tse_ddr_clock_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_sgdma_tx_m_read_to_tse_ddr_clock_bridge_s1_module;

                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal internal_tse_ddr_clock_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_sgdma_rx_m_write_granted_slave_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_tx_m_read_granted_slave_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal module_input37 :  STD_LOGIC;
                signal module_input38 :  STD_LOGIC;
                signal module_input39 :  STD_LOGIC;
                signal sgdma_rx_m_write_arbiterlock :  STD_LOGIC;
                signal sgdma_rx_m_write_arbiterlock2 :  STD_LOGIC;
                signal sgdma_rx_m_write_continuerequest :  STD_LOGIC;
                signal sgdma_rx_m_write_saved_grant_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_arbiterlock :  STD_LOGIC;
                signal sgdma_tx_m_read_arbiterlock2 :  STD_LOGIC;
                signal sgdma_tx_m_read_continuerequest :  STD_LOGIC;
                signal sgdma_tx_m_read_rdv_fifo_empty_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_rdv_fifo_output_from_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_saved_grant_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal shifted_address_to_tse_ddr_clock_bridge_s1_from_sgdma_rx_m_write :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_tse_ddr_clock_bridge_s1_from_sgdma_tx_m_read :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_allgrants :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_any_continuerequest :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_arb_counter_enable :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_arb_share_counter :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_arb_share_set_values :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_begins_xfer :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_end_xfer :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_firsttransfer :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_in_a_read_cycle :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_in_a_write_cycle :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_non_bursting_master_requests :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_reg_firsttransfer :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_slavearbiterlockenable :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_unreg_firsttransfer :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_waits_for_read :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_tse_ddr_clock_bridge_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT tse_ddr_clock_bridge_s1_end_xfer;
    end if;

  end process;

  tse_ddr_clock_bridge_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 OR internal_sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1));
  --assign tse_ddr_clock_bridge_s1_readdata_from_sa = tse_ddr_clock_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  tse_ddr_clock_bridge_s1_readdata_from_sa <= tse_ddr_clock_bridge_s1_readdata;
  internal_sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_rx_m_write_address_to_slave(31 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (sgdma_rx_m_write_write))) AND sgdma_rx_m_write_write;
  --assign tse_ddr_clock_bridge_s1_waitrequest_from_sa = tse_ddr_clock_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_tse_ddr_clock_bridge_s1_waitrequest_from_sa <= tse_ddr_clock_bridge_s1_waitrequest;
  --tse_ddr_clock_bridge_s1_arb_share_counter set values, which is an e_mux
  tse_ddr_clock_bridge_s1_arb_share_set_values <= std_logic'('1');
  --tse_ddr_clock_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  tse_ddr_clock_bridge_s1_non_bursting_master_requests <= ((internal_sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 OR internal_sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1) OR internal_sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1) OR internal_sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1;
  --tse_ddr_clock_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  tse_ddr_clock_bridge_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --tse_ddr_clock_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  tse_ddr_clock_bridge_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(tse_ddr_clock_bridge_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_ddr_clock_bridge_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(tse_ddr_clock_bridge_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_ddr_clock_bridge_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --tse_ddr_clock_bridge_s1_allgrants all slave grants, which is an e_mux
  tse_ddr_clock_bridge_s1_allgrants <= (((or_reduce(tse_ddr_clock_bridge_s1_grant_vector)) OR (or_reduce(tse_ddr_clock_bridge_s1_grant_vector))) OR (or_reduce(tse_ddr_clock_bridge_s1_grant_vector))) OR (or_reduce(tse_ddr_clock_bridge_s1_grant_vector));
  --tse_ddr_clock_bridge_s1_end_xfer assignment, which is an e_assign
  tse_ddr_clock_bridge_s1_end_xfer <= NOT ((tse_ddr_clock_bridge_s1_waits_for_read OR tse_ddr_clock_bridge_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_tse_ddr_clock_bridge_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_tse_ddr_clock_bridge_s1 <= tse_ddr_clock_bridge_s1_end_xfer AND (((NOT tse_ddr_clock_bridge_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --tse_ddr_clock_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  tse_ddr_clock_bridge_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_tse_ddr_clock_bridge_s1 AND tse_ddr_clock_bridge_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_tse_ddr_clock_bridge_s1 AND NOT tse_ddr_clock_bridge_s1_non_bursting_master_requests));
  --tse_ddr_clock_bridge_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_ddr_clock_bridge_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(tse_ddr_clock_bridge_s1_arb_counter_enable) = '1' then 
        tse_ddr_clock_bridge_s1_arb_share_counter <= tse_ddr_clock_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --tse_ddr_clock_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_ddr_clock_bridge_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(tse_ddr_clock_bridge_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_tse_ddr_clock_bridge_s1)) OR ((end_xfer_arb_share_counter_term_tse_ddr_clock_bridge_s1 AND NOT tse_ddr_clock_bridge_s1_non_bursting_master_requests)))) = '1' then 
        tse_ddr_clock_bridge_s1_slavearbiterlockenable <= tse_ddr_clock_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sgdma_rx/m_write tse_ddr_clock_bridge/s1 arbiterlock, which is an e_assign
  sgdma_rx_m_write_arbiterlock <= tse_ddr_clock_bridge_s1_slavearbiterlockenable AND sgdma_rx_m_write_continuerequest;
  --tse_ddr_clock_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  tse_ddr_clock_bridge_s1_slavearbiterlockenable2 <= tse_ddr_clock_bridge_s1_arb_share_counter_next_value;
  --sgdma_rx/m_write tse_ddr_clock_bridge/s1 arbiterlock2, which is an e_assign
  sgdma_rx_m_write_arbiterlock2 <= tse_ddr_clock_bridge_s1_slavearbiterlockenable2 AND sgdma_rx_m_write_continuerequest;
  --sgdma_tx/m_read tse_ddr_clock_bridge/s1 arbiterlock, which is an e_assign
  sgdma_tx_m_read_arbiterlock <= tse_ddr_clock_bridge_s1_slavearbiterlockenable AND sgdma_tx_m_read_continuerequest;
  --sgdma_tx/m_read tse_ddr_clock_bridge/s1 arbiterlock2, which is an e_assign
  sgdma_tx_m_read_arbiterlock2 <= tse_ddr_clock_bridge_s1_slavearbiterlockenable2 AND sgdma_tx_m_read_continuerequest;
  --sgdma_tx/m_read granted tse_ddr_clock_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_tx_m_read_granted_slave_tse_ddr_clock_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_tx_m_read_granted_slave_tse_ddr_clock_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_tx_m_read_saved_grant_tse_ddr_clock_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((tse_ddr_clock_bridge_s1_arbitration_holdoff_internal OR NOT internal_sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_tx_m_read_granted_slave_tse_ddr_clock_bridge_s1))))));
    end if;

  end process;

  --sgdma_tx_m_read_continuerequest continued request, which is an e_mux
  sgdma_tx_m_read_continuerequest <= last_cycle_sgdma_tx_m_read_granted_slave_tse_ddr_clock_bridge_s1 AND internal_sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1;
  --tse_ddr_clock_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  tse_ddr_clock_bridge_s1_any_continuerequest <= sgdma_tx_m_read_continuerequest OR sgdma_rx_m_write_continuerequest;
  internal_sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 <= internal_sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 AND NOT (sgdma_tx_m_read_arbiterlock);
  --tse_ddr_clock_bridge_s1_writedata mux, which is an e_mux
  tse_ddr_clock_bridge_s1_writedata <= sgdma_rx_m_write_writedata;
  --assign tse_ddr_clock_bridge_s1_endofpacket_from_sa = tse_ddr_clock_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  tse_ddr_clock_bridge_s1_endofpacket_from_sa <= tse_ddr_clock_bridge_s1_endofpacket;
  internal_sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_tx_m_read_address_to_slave(31 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000000000000000000000000000000")))) AND (sgdma_tx_m_read_read))) AND sgdma_tx_m_read_read;
  --assign tse_ddr_clock_bridge_s1_readdatavalid_from_sa = tse_ddr_clock_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  tse_ddr_clock_bridge_s1_readdatavalid_from_sa <= tse_ddr_clock_bridge_s1_readdatavalid;
  --sgdma_rx/m_write granted tse_ddr_clock_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_rx_m_write_granted_slave_tse_ddr_clock_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_rx_m_write_granted_slave_tse_ddr_clock_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_rx_m_write_saved_grant_tse_ddr_clock_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((tse_ddr_clock_bridge_s1_arbitration_holdoff_internal OR NOT internal_sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_rx_m_write_granted_slave_tse_ddr_clock_bridge_s1))))));
    end if;

  end process;

  --sgdma_rx_m_write_continuerequest continued request, which is an e_mux
  sgdma_rx_m_write_continuerequest <= last_cycle_sgdma_rx_m_write_granted_slave_tse_ddr_clock_bridge_s1 AND internal_sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1;
  internal_sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 <= internal_sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 AND NOT ((((sgdma_tx_m_read_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_tx_m_read_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_tx_m_read_latency_counter)))))))))) OR sgdma_rx_m_write_arbiterlock));
  --unique name for tse_ddr_clock_bridge_s1_move_on_to_next_transaction, which is an e_assign
  tse_ddr_clock_bridge_s1_move_on_to_next_transaction <= tse_ddr_clock_bridge_s1_readdatavalid_from_sa;
  --rdv_fifo_for_sgdma_tx_m_read_to_tse_ddr_clock_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_sgdma_tx_m_read_to_tse_ddr_clock_bridge_s1 : rdv_fifo_for_sgdma_tx_m_read_to_tse_ddr_clock_bridge_s1_module
    port map(
      data_out => sgdma_tx_m_read_rdv_fifo_output_from_tse_ddr_clock_bridge_s1,
      empty => open,
      fifo_contains_ones_n => sgdma_tx_m_read_rdv_fifo_empty_tse_ddr_clock_bridge_s1,
      full => open,
      clear_fifo => module_input37,
      clk => clk,
      data_in => internal_sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1,
      read => tse_ddr_clock_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input38,
      write => module_input39
    );

  module_input37 <= std_logic'('0');
  module_input38 <= std_logic'('0');
  module_input39 <= in_a_read_cycle AND NOT tse_ddr_clock_bridge_s1_waits_for_read;

  sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1_shift_register <= NOT sgdma_tx_m_read_rdv_fifo_empty_tse_ddr_clock_bridge_s1;
  --local readdatavalid sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1, which is an e_mux
  sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1 <= ((tse_ddr_clock_bridge_s1_readdatavalid_from_sa AND sgdma_tx_m_read_rdv_fifo_output_from_tse_ddr_clock_bridge_s1)) AND NOT sgdma_tx_m_read_rdv_fifo_empty_tse_ddr_clock_bridge_s1;
  --allow new arb cycle for tse_ddr_clock_bridge/s1, which is an e_assign
  tse_ddr_clock_bridge_s1_allow_new_arb_cycle <= NOT sgdma_rx_m_write_arbiterlock AND NOT sgdma_tx_m_read_arbiterlock;
  --sgdma_tx/m_read assignment into master qualified-requests vector for tse_ddr_clock_bridge/s1, which is an e_assign
  tse_ddr_clock_bridge_s1_master_qreq_vector(0) <= internal_sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1;
  --sgdma_tx/m_read grant tse_ddr_clock_bridge/s1, which is an e_assign
  internal_sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 <= tse_ddr_clock_bridge_s1_grant_vector(0);
  --sgdma_tx/m_read saved-grant tse_ddr_clock_bridge/s1, which is an e_assign
  sgdma_tx_m_read_saved_grant_tse_ddr_clock_bridge_s1 <= tse_ddr_clock_bridge_s1_arb_winner(0) AND internal_sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1;
  --sgdma_rx/m_write assignment into master qualified-requests vector for tse_ddr_clock_bridge/s1, which is an e_assign
  tse_ddr_clock_bridge_s1_master_qreq_vector(1) <= internal_sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1;
  --sgdma_rx/m_write grant tse_ddr_clock_bridge/s1, which is an e_assign
  internal_sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 <= tse_ddr_clock_bridge_s1_grant_vector(1);
  --sgdma_rx/m_write saved-grant tse_ddr_clock_bridge/s1, which is an e_assign
  sgdma_rx_m_write_saved_grant_tse_ddr_clock_bridge_s1 <= tse_ddr_clock_bridge_s1_arb_winner(1) AND internal_sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1;
  --tse_ddr_clock_bridge/s1 chosen-master double-vector, which is an e_assign
  tse_ddr_clock_bridge_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((tse_ddr_clock_bridge_s1_master_qreq_vector & tse_ddr_clock_bridge_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT tse_ddr_clock_bridge_s1_master_qreq_vector & NOT tse_ddr_clock_bridge_s1_master_qreq_vector))) + (std_logic_vector'("000") & (tse_ddr_clock_bridge_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  tse_ddr_clock_bridge_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((tse_ddr_clock_bridge_s1_allow_new_arb_cycle AND or_reduce(tse_ddr_clock_bridge_s1_grant_vector)))) = '1'), tse_ddr_clock_bridge_s1_grant_vector, tse_ddr_clock_bridge_s1_saved_chosen_master_vector);
  --saved tse_ddr_clock_bridge_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_ddr_clock_bridge_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(tse_ddr_clock_bridge_s1_allow_new_arb_cycle) = '1' then 
        tse_ddr_clock_bridge_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(tse_ddr_clock_bridge_s1_grant_vector)) = '1'), tse_ddr_clock_bridge_s1_grant_vector, tse_ddr_clock_bridge_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  tse_ddr_clock_bridge_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((tse_ddr_clock_bridge_s1_chosen_master_double_vector(1) OR tse_ddr_clock_bridge_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((tse_ddr_clock_bridge_s1_chosen_master_double_vector(0) OR tse_ddr_clock_bridge_s1_chosen_master_double_vector(2)))));
  --tse_ddr_clock_bridge/s1 chosen master rotated left, which is an e_assign
  tse_ddr_clock_bridge_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(tse_ddr_clock_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(tse_ddr_clock_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --tse_ddr_clock_bridge/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_ddr_clock_bridge_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(tse_ddr_clock_bridge_s1_grant_vector)) = '1' then 
        tse_ddr_clock_bridge_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(tse_ddr_clock_bridge_s1_end_xfer) = '1'), tse_ddr_clock_bridge_s1_chosen_master_rot_left, tse_ddr_clock_bridge_s1_grant_vector);
      end if;
    end if;

  end process;

  --tse_ddr_clock_bridge_s1_reset_n assignment, which is an e_assign
  tse_ddr_clock_bridge_s1_reset_n <= reset_n;
  --tse_ddr_clock_bridge_s1_firsttransfer first transaction, which is an e_assign
  tse_ddr_clock_bridge_s1_firsttransfer <= A_WE_StdLogic((std_logic'(tse_ddr_clock_bridge_s1_begins_xfer) = '1'), tse_ddr_clock_bridge_s1_unreg_firsttransfer, tse_ddr_clock_bridge_s1_reg_firsttransfer);
  --tse_ddr_clock_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  tse_ddr_clock_bridge_s1_unreg_firsttransfer <= NOT ((tse_ddr_clock_bridge_s1_slavearbiterlockenable AND tse_ddr_clock_bridge_s1_any_continuerequest));
  --tse_ddr_clock_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_ddr_clock_bridge_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(tse_ddr_clock_bridge_s1_begins_xfer) = '1' then 
        tse_ddr_clock_bridge_s1_reg_firsttransfer <= tse_ddr_clock_bridge_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --tse_ddr_clock_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  tse_ddr_clock_bridge_s1_beginbursttransfer_internal <= tse_ddr_clock_bridge_s1_begins_xfer;
  --tse_ddr_clock_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  tse_ddr_clock_bridge_s1_arbitration_holdoff_internal <= tse_ddr_clock_bridge_s1_begins_xfer AND tse_ddr_clock_bridge_s1_firsttransfer;
  --tse_ddr_clock_bridge_s1_read assignment, which is an e_mux
  tse_ddr_clock_bridge_s1_read <= internal_sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 AND sgdma_tx_m_read_read;
  --tse_ddr_clock_bridge_s1_write assignment, which is an e_mux
  tse_ddr_clock_bridge_s1_write <= internal_sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 AND sgdma_rx_m_write_write;
  shifted_address_to_tse_ddr_clock_bridge_s1_from_sgdma_rx_m_write <= sgdma_rx_m_write_address_to_slave;
  --tse_ddr_clock_bridge_s1_address mux, which is an e_mux
  tse_ddr_clock_bridge_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1)) = '1'), (A_SRL(shifted_address_to_tse_ddr_clock_bridge_s1_from_sgdma_rx_m_write,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_tse_ddr_clock_bridge_s1_from_sgdma_tx_m_read,std_logic_vector'("00000000000000000000000000000010")))), 23);
  shifted_address_to_tse_ddr_clock_bridge_s1_from_sgdma_tx_m_read <= sgdma_tx_m_read_address_to_slave;
  --slaveid tse_ddr_clock_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  tse_ddr_clock_bridge_s1_nativeaddress <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1)) = '1'), (A_SRL(sgdma_rx_m_write_address_to_slave,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(sgdma_tx_m_read_address_to_slave,std_logic_vector'("00000000000000000000000000000010")))), 23);
  --d1_tse_ddr_clock_bridge_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_tse_ddr_clock_bridge_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_tse_ddr_clock_bridge_s1_end_xfer <= tse_ddr_clock_bridge_s1_end_xfer;
    end if;

  end process;

  --tse_ddr_clock_bridge_s1_waits_for_read in a cycle, which is an e_mux
  tse_ddr_clock_bridge_s1_waits_for_read <= tse_ddr_clock_bridge_s1_in_a_read_cycle AND internal_tse_ddr_clock_bridge_s1_waitrequest_from_sa;
  --tse_ddr_clock_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  tse_ddr_clock_bridge_s1_in_a_read_cycle <= internal_sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 AND sgdma_tx_m_read_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= tse_ddr_clock_bridge_s1_in_a_read_cycle;
  --tse_ddr_clock_bridge_s1_waits_for_write in a cycle, which is an e_mux
  tse_ddr_clock_bridge_s1_waits_for_write <= tse_ddr_clock_bridge_s1_in_a_write_cycle AND internal_tse_ddr_clock_bridge_s1_waitrequest_from_sa;
  --tse_ddr_clock_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  tse_ddr_clock_bridge_s1_in_a_write_cycle <= internal_sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 AND sgdma_rx_m_write_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= tse_ddr_clock_bridge_s1_in_a_write_cycle;
  wait_for_tse_ddr_clock_bridge_s1_counter <= std_logic'('0');
  --tse_ddr_clock_bridge_s1_byteenable byte enable port mux, which is an e_mux
  tse_ddr_clock_bridge_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (sgdma_rx_m_write_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 <= internal_sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 <= internal_sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 <= internal_sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 <= internal_sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 <= internal_sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 <= internal_sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1;
  --vhdl renameroo for output signals
  tse_ddr_clock_bridge_s1_waitrequest_from_sa <= internal_tse_ddr_clock_bridge_s1_waitrequest_from_sa;
--synthesis translate_off
    --tse_ddr_clock_bridge/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line56 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line56, now);
          write(write_line56, string'(": "));
          write(write_line56, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line56.all);
          deallocate (write_line56);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line57 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(sgdma_rx_m_write_saved_grant_tse_ddr_clock_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(sgdma_tx_m_read_saved_grant_tse_ddr_clock_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line57, now);
          write(write_line57, string'(": "));
          write(write_line57, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line57.all);
          deallocate (write_line57);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_module;


architecture europa of selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_17 :  STD_LOGIC;
                signal full_18 :  STD_LOGIC;
                signal full_19 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_20 :  STD_LOGIC;
                signal full_21 :  STD_LOGIC;
                signal full_22 :  STD_LOGIC;
                signal full_23 :  STD_LOGIC;
                signal full_24 :  STD_LOGIC;
                signal full_25 :  STD_LOGIC;
                signal full_26 :  STD_LOGIC;
                signal full_27 :  STD_LOGIC;
                signal full_28 :  STD_LOGIC;
                signal full_29 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_30 :  STD_LOGIC;
                signal full_31 :  STD_LOGIC;
                signal full_32 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p16_full_16 :  STD_LOGIC;
                signal p16_stage_16 :  STD_LOGIC;
                signal p17_full_17 :  STD_LOGIC;
                signal p17_stage_17 :  STD_LOGIC;
                signal p18_full_18 :  STD_LOGIC;
                signal p18_stage_18 :  STD_LOGIC;
                signal p19_full_19 :  STD_LOGIC;
                signal p19_stage_19 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p20_full_20 :  STD_LOGIC;
                signal p20_stage_20 :  STD_LOGIC;
                signal p21_full_21 :  STD_LOGIC;
                signal p21_stage_21 :  STD_LOGIC;
                signal p22_full_22 :  STD_LOGIC;
                signal p22_stage_22 :  STD_LOGIC;
                signal p23_full_23 :  STD_LOGIC;
                signal p23_stage_23 :  STD_LOGIC;
                signal p24_full_24 :  STD_LOGIC;
                signal p24_stage_24 :  STD_LOGIC;
                signal p25_full_25 :  STD_LOGIC;
                signal p25_stage_25 :  STD_LOGIC;
                signal p26_full_26 :  STD_LOGIC;
                signal p26_stage_26 :  STD_LOGIC;
                signal p27_full_27 :  STD_LOGIC;
                signal p27_stage_27 :  STD_LOGIC;
                signal p28_full_28 :  STD_LOGIC;
                signal p28_stage_28 :  STD_LOGIC;
                signal p29_full_29 :  STD_LOGIC;
                signal p29_stage_29 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p30_full_30 :  STD_LOGIC;
                signal p30_stage_30 :  STD_LOGIC;
                signal p31_full_31 :  STD_LOGIC;
                signal p31_stage_31 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_16 :  STD_LOGIC;
                signal stage_17 :  STD_LOGIC;
                signal stage_18 :  STD_LOGIC;
                signal stage_19 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_20 :  STD_LOGIC;
                signal stage_21 :  STD_LOGIC;
                signal stage_22 :  STD_LOGIC;
                signal stage_23 :  STD_LOGIC;
                signal stage_24 :  STD_LOGIC;
                signal stage_25 :  STD_LOGIC;
                signal stage_26 :  STD_LOGIC;
                signal stage_27 :  STD_LOGIC;
                signal stage_28 :  STD_LOGIC;
                signal stage_29 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_30 :  STD_LOGIC;
                signal stage_31 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (6 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_31;
  empty <= NOT(full_0);
  full_32 <= std_logic'('0');
  --data_31, which is an e_mux
  p31_stage_31 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_32 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_31))))) = '1' then 
        if std_logic'(((sync_reset AND full_31) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_32))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_31 <= std_logic'('0');
        else
          stage_31 <= p31_stage_31;
        end if;
      end if;
    end if;

  end process;

  --control_31, which is an e_mux
  p31_full_31 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_31, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_31 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_31 <= std_logic'('0');
        else
          full_31 <= p31_full_31;
        end if;
      end if;
    end if;

  end process;

  --data_30, which is an e_mux
  p30_stage_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_31 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_31);
  --data_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_30))))) = '1' then 
        if std_logic'(((sync_reset AND full_30) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_31))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_30 <= std_logic'('0');
        else
          stage_30 <= p30_stage_30;
        end if;
      end if;
    end if;

  end process;

  --control_30, which is an e_mux
  p30_full_30 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_29, full_31);
  --control_reg_30, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_30 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_30 <= std_logic'('0');
        else
          full_30 <= p30_full_30;
        end if;
      end if;
    end if;

  end process;

  --data_29, which is an e_mux
  p29_stage_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_30 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_30);
  --data_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_29))))) = '1' then 
        if std_logic'(((sync_reset AND full_29) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_30))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_29 <= std_logic'('0');
        else
          stage_29 <= p29_stage_29;
        end if;
      end if;
    end if;

  end process;

  --control_29, which is an e_mux
  p29_full_29 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_28, full_30);
  --control_reg_29, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_29 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_29 <= std_logic'('0');
        else
          full_29 <= p29_full_29;
        end if;
      end if;
    end if;

  end process;

  --data_28, which is an e_mux
  p28_stage_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_29 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_29);
  --data_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_28))))) = '1' then 
        if std_logic'(((sync_reset AND full_28) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_29))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_28 <= std_logic'('0');
        else
          stage_28 <= p28_stage_28;
        end if;
      end if;
    end if;

  end process;

  --control_28, which is an e_mux
  p28_full_28 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_27, full_29);
  --control_reg_28, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_28 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_28 <= std_logic'('0');
        else
          full_28 <= p28_full_28;
        end if;
      end if;
    end if;

  end process;

  --data_27, which is an e_mux
  p27_stage_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_28 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_28);
  --data_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_27))))) = '1' then 
        if std_logic'(((sync_reset AND full_27) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_28))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_27 <= std_logic'('0');
        else
          stage_27 <= p27_stage_27;
        end if;
      end if;
    end if;

  end process;

  --control_27, which is an e_mux
  p27_full_27 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_26, full_28);
  --control_reg_27, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_27 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_27 <= std_logic'('0');
        else
          full_27 <= p27_full_27;
        end if;
      end if;
    end if;

  end process;

  --data_26, which is an e_mux
  p26_stage_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_27 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_27);
  --data_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_26))))) = '1' then 
        if std_logic'(((sync_reset AND full_26) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_27))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_26 <= std_logic'('0');
        else
          stage_26 <= p26_stage_26;
        end if;
      end if;
    end if;

  end process;

  --control_26, which is an e_mux
  p26_full_26 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_25, full_27);
  --control_reg_26, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_26 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_26 <= std_logic'('0');
        else
          full_26 <= p26_full_26;
        end if;
      end if;
    end if;

  end process;

  --data_25, which is an e_mux
  p25_stage_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_26 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_26);
  --data_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_25))))) = '1' then 
        if std_logic'(((sync_reset AND full_25) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_26))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_25 <= std_logic'('0');
        else
          stage_25 <= p25_stage_25;
        end if;
      end if;
    end if;

  end process;

  --control_25, which is an e_mux
  p25_full_25 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_24, full_26);
  --control_reg_25, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_25 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_25 <= std_logic'('0');
        else
          full_25 <= p25_full_25;
        end if;
      end if;
    end if;

  end process;

  --data_24, which is an e_mux
  p24_stage_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_25 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_25);
  --data_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_24))))) = '1' then 
        if std_logic'(((sync_reset AND full_24) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_25))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_24 <= std_logic'('0');
        else
          stage_24 <= p24_stage_24;
        end if;
      end if;
    end if;

  end process;

  --control_24, which is an e_mux
  p24_full_24 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_23, full_25);
  --control_reg_24, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_24 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_24 <= std_logic'('0');
        else
          full_24 <= p24_full_24;
        end if;
      end if;
    end if;

  end process;

  --data_23, which is an e_mux
  p23_stage_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_24 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_24);
  --data_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_23))))) = '1' then 
        if std_logic'(((sync_reset AND full_23) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_24))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_23 <= std_logic'('0');
        else
          stage_23 <= p23_stage_23;
        end if;
      end if;
    end if;

  end process;

  --control_23, which is an e_mux
  p23_full_23 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_22, full_24);
  --control_reg_23, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_23 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_23 <= std_logic'('0');
        else
          full_23 <= p23_full_23;
        end if;
      end if;
    end if;

  end process;

  --data_22, which is an e_mux
  p22_stage_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_23 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_23);
  --data_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_22))))) = '1' then 
        if std_logic'(((sync_reset AND full_22) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_23))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_22 <= std_logic'('0');
        else
          stage_22 <= p22_stage_22;
        end if;
      end if;
    end if;

  end process;

  --control_22, which is an e_mux
  p22_full_22 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_21, full_23);
  --control_reg_22, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_22 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_22 <= std_logic'('0');
        else
          full_22 <= p22_full_22;
        end if;
      end if;
    end if;

  end process;

  --data_21, which is an e_mux
  p21_stage_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_22 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_22);
  --data_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_21))))) = '1' then 
        if std_logic'(((sync_reset AND full_21) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_22))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_21 <= std_logic'('0');
        else
          stage_21 <= p21_stage_21;
        end if;
      end if;
    end if;

  end process;

  --control_21, which is an e_mux
  p21_full_21 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_20, full_22);
  --control_reg_21, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_21 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_21 <= std_logic'('0');
        else
          full_21 <= p21_full_21;
        end if;
      end if;
    end if;

  end process;

  --data_20, which is an e_mux
  p20_stage_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_21 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_21);
  --data_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_20))))) = '1' then 
        if std_logic'(((sync_reset AND full_20) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_21))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_20 <= std_logic'('0');
        else
          stage_20 <= p20_stage_20;
        end if;
      end if;
    end if;

  end process;

  --control_20, which is an e_mux
  p20_full_20 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_19, full_21);
  --control_reg_20, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_20 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_20 <= std_logic'('0');
        else
          full_20 <= p20_full_20;
        end if;
      end if;
    end if;

  end process;

  --data_19, which is an e_mux
  p19_stage_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_20 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_20);
  --data_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_19))))) = '1' then 
        if std_logic'(((sync_reset AND full_19) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_20))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_19 <= std_logic'('0');
        else
          stage_19 <= p19_stage_19;
        end if;
      end if;
    end if;

  end process;

  --control_19, which is an e_mux
  p19_full_19 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_18, full_20);
  --control_reg_19, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_19 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_19 <= std_logic'('0');
        else
          full_19 <= p19_full_19;
        end if;
      end if;
    end if;

  end process;

  --data_18, which is an e_mux
  p18_stage_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_19 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_19);
  --data_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_18))))) = '1' then 
        if std_logic'(((sync_reset AND full_18) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_19))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_18 <= std_logic'('0');
        else
          stage_18 <= p18_stage_18;
        end if;
      end if;
    end if;

  end process;

  --control_18, which is an e_mux
  p18_full_18 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_17, full_19);
  --control_reg_18, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_18 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_18 <= std_logic'('0');
        else
          full_18 <= p18_full_18;
        end if;
      end if;
    end if;

  end process;

  --data_17, which is an e_mux
  p17_stage_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_18 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_18);
  --data_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_17))))) = '1' then 
        if std_logic'(((sync_reset AND full_17) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_18))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_17 <= std_logic'('0');
        else
          stage_17 <= p17_stage_17;
        end if;
      end if;
    end if;

  end process;

  --control_17, which is an e_mux
  p17_full_17 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_16, full_18);
  --control_reg_17, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_17 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_17 <= std_logic'('0');
        else
          full_17 <= p17_full_17;
        end if;
      end if;
    end if;

  end process;

  --data_16, which is an e_mux
  p16_stage_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_17 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_17);
  --data_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_16))))) = '1' then 
        if std_logic'(((sync_reset AND full_16) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_17))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_16 <= std_logic'('0');
        else
          stage_16 <= p16_stage_16;
        end if;
      end if;
    end if;

  end process;

  --control_16, which is an e_mux
  p16_full_16 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_15, full_17);
  --control_reg_16, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_16 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_16 <= std_logic'('0');
        else
          full_16 <= p16_full_16;
        end if;
      end if;
    end if;

  end process;

  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_16);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_14, full_16);
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 7);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 7);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 7);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity tse_ddr_clock_bridge_m1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                 signal sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal tse_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal tse_ddr_clock_bridge_m1_granted_sdram_s1 : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1 : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_requests_sdram_s1 : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal tse_ddr_clock_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal tse_ddr_clock_bridge_m1_latency_counter : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_ddr_clock_bridge_m1_readdatavalid : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_reset_n : OUT STD_LOGIC;
                 signal tse_ddr_clock_bridge_m1_waitrequest : OUT STD_LOGIC
              );
end entity tse_ddr_clock_bridge_m1_arbitrator;


architecture europa of tse_ddr_clock_bridge_m1_arbitrator is
component selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_module;

                signal active_and_waiting_last_time :  STD_LOGIC;
                signal empty_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo :  STD_LOGIC;
                signal full_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo :  STD_LOGIC;
                signal internal_tse_ddr_clock_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_tse_ddr_clock_bridge_m1_latency_counter :  STD_LOGIC;
                signal internal_tse_ddr_clock_bridge_m1_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal module_input40 :  STD_LOGIC;
                signal module_input41 :  STD_LOGIC;
                signal module_input42 :  STD_LOGIC;
                signal p1_tse_ddr_clock_bridge_m1_latency_counter :  STD_LOGIC;
                signal pre_flush_tse_ddr_clock_bridge_m1_readdatavalid :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal read_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo :  STD_LOGIC;
                signal sdram_s1_readdata_from_sa_part_selected_by_negative_dbs :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_output :  STD_LOGIC;
                signal selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_output_sdram_s1 :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal tse_ddr_clock_bridge_m1_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tse_ddr_clock_bridge_m1_is_granted_some_slave :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_read_but_no_slave_selected :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_read_last_time :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_run :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_write_last_time :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal write_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 OR NOT tse_ddr_clock_bridge_m1_requests_sdram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((tse_ddr_clock_bridge_m1_granted_sdram_s1 OR NOT tse_ddr_clock_bridge_m1_qualified_request_sdram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 OR NOT ((tse_ddr_clock_bridge_m1_read OR tse_ddr_clock_bridge_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((tse_ddr_clock_bridge_m1_read OR tse_ddr_clock_bridge_m1_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 OR NOT ((tse_ddr_clock_bridge_m1_read OR tse_ddr_clock_bridge_m1_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((tse_ddr_clock_bridge_m1_read OR tse_ddr_clock_bridge_m1_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  tse_ddr_clock_bridge_m1_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_tse_ddr_clock_bridge_m1_address_to_slave <= tse_ddr_clock_bridge_m1_address(24 DOWNTO 0);
  --tse_ddr_clock_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_ddr_clock_bridge_m1_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      tse_ddr_clock_bridge_m1_read_but_no_slave_selected <= (tse_ddr_clock_bridge_m1_read AND tse_ddr_clock_bridge_m1_run) AND NOT tse_ddr_clock_bridge_m1_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  tse_ddr_clock_bridge_m1_is_granted_some_slave <= tse_ddr_clock_bridge_m1_granted_sdram_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_tse_ddr_clock_bridge_m1_readdatavalid <= tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  tse_ddr_clock_bridge_m1_readdatavalid <= tse_ddr_clock_bridge_m1_read_but_no_slave_selected OR pre_flush_tse_ddr_clock_bridge_m1_readdatavalid;
  --Negative Dynamic Bus-sizing mux.
  --this mux selects the correct half of the 
  --wide data coming from the slave sdram/s1 
  sdram_s1_readdata_from_sa_part_selected_by_negative_dbs <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_output_sdram_s1))) = std_logic_vector'("00000000000000000000000000000000"))), sdram_s1_readdata_from_sa(31 DOWNTO 0), sdram_s1_readdata_from_sa(63 DOWNTO 32));
  --read_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo fifo read, which is an e_mux
  read_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo <= tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1;
  --write_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo fifo write, which is an e_mux
  write_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo <= (tse_ddr_clock_bridge_m1_read AND tse_ddr_clock_bridge_m1_run) AND tse_ddr_clock_bridge_m1_requests_sdram_s1;
  selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_output_sdram_s1 <= selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_output;
  --selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo, which is an e_fifo_with_registered_outputs
  selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo : selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_module
    port map(
      data_out => selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo_output,
      empty => empty_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo,
      fifo_contains_ones_n => open,
      full => full_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo,
      clear_fifo => module_input40,
      clk => clk,
      data_in => module_input41,
      read => read_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo,
      reset_n => reset_n,
      sync_reset => module_input42,
      write => write_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo
    );

  module_input40 <= std_logic'('0');
  module_input41 <= internal_tse_ddr_clock_bridge_m1_address_to_slave(2);
  module_input42 <= std_logic'('0');

  --tse_ddr_clock_bridge/m1 readdata mux, which is an e_mux
  tse_ddr_clock_bridge_m1_readdata <= sdram_s1_readdata_from_sa_part_selected_by_negative_dbs;
  --actual waitrequest port, which is an e_assign
  internal_tse_ddr_clock_bridge_m1_waitrequest <= NOT tse_ddr_clock_bridge_m1_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_tse_ddr_clock_bridge_m1_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_tse_ddr_clock_bridge_m1_latency_counter <= p1_tse_ddr_clock_bridge_m1_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_tse_ddr_clock_bridge_m1_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((tse_ddr_clock_bridge_m1_run AND tse_ddr_clock_bridge_m1_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_tse_ddr_clock_bridge_m1_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_tse_ddr_clock_bridge_m1_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --tse_ddr_clock_bridge_m1_reset_n assignment, which is an e_assign
  tse_ddr_clock_bridge_m1_reset_n <= reset_n;
  --vhdl renameroo for output signals
  tse_ddr_clock_bridge_m1_address_to_slave <= internal_tse_ddr_clock_bridge_m1_address_to_slave;
  --vhdl renameroo for output signals
  tse_ddr_clock_bridge_m1_latency_counter <= internal_tse_ddr_clock_bridge_m1_latency_counter;
  --vhdl renameroo for output signals
  tse_ddr_clock_bridge_m1_waitrequest <= internal_tse_ddr_clock_bridge_m1_waitrequest;
--synthesis translate_off
    --tse_ddr_clock_bridge_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        tse_ddr_clock_bridge_m1_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        tse_ddr_clock_bridge_m1_address_last_time <= tse_ddr_clock_bridge_m1_address;
      end if;

    end process;

    --tse_ddr_clock_bridge/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_tse_ddr_clock_bridge_m1_waitrequest AND ((tse_ddr_clock_bridge_m1_read OR tse_ddr_clock_bridge_m1_write));
      end if;

    end process;

    --tse_ddr_clock_bridge_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line58 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((tse_ddr_clock_bridge_m1_address /= tse_ddr_clock_bridge_m1_address_last_time))))) = '1' then 
          write(write_line58, now);
          write(write_line58, string'(": "));
          write(write_line58, string'("tse_ddr_clock_bridge_m1_address did not heed wait!!!"));
          write(output, write_line58.all);
          deallocate (write_line58);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --tse_ddr_clock_bridge_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        tse_ddr_clock_bridge_m1_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        tse_ddr_clock_bridge_m1_byteenable_last_time <= tse_ddr_clock_bridge_m1_byteenable;
      end if;

    end process;

    --tse_ddr_clock_bridge_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line59 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((tse_ddr_clock_bridge_m1_byteenable /= tse_ddr_clock_bridge_m1_byteenable_last_time))))) = '1' then 
          write(write_line59, now);
          write(write_line59, string'(": "));
          write(write_line59, string'("tse_ddr_clock_bridge_m1_byteenable did not heed wait!!!"));
          write(output, write_line59.all);
          deallocate (write_line59);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --tse_ddr_clock_bridge_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        tse_ddr_clock_bridge_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        tse_ddr_clock_bridge_m1_read_last_time <= tse_ddr_clock_bridge_m1_read;
      end if;

    end process;

    --tse_ddr_clock_bridge_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line60 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(tse_ddr_clock_bridge_m1_read) /= std_logic'(tse_ddr_clock_bridge_m1_read_last_time)))))) = '1' then 
          write(write_line60, now);
          write(write_line60, string'(": "));
          write(write_line60, string'("tse_ddr_clock_bridge_m1_read did not heed wait!!!"));
          write(output, write_line60.all);
          deallocate (write_line60);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --tse_ddr_clock_bridge_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        tse_ddr_clock_bridge_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        tse_ddr_clock_bridge_m1_write_last_time <= tse_ddr_clock_bridge_m1_write;
      end if;

    end process;

    --tse_ddr_clock_bridge_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line61 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(tse_ddr_clock_bridge_m1_write) /= std_logic'(tse_ddr_clock_bridge_m1_write_last_time)))))) = '1' then 
          write(write_line61, now);
          write(write_line61, string'(": "));
          write(write_line61, string'("tse_ddr_clock_bridge_m1_write did not heed wait!!!"));
          write(output, write_line61.all);
          deallocate (write_line61);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --tse_ddr_clock_bridge_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        tse_ddr_clock_bridge_m1_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        tse_ddr_clock_bridge_m1_writedata_last_time <= tse_ddr_clock_bridge_m1_writedata;
      end if;

    end process;

    --tse_ddr_clock_bridge_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line62 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((tse_ddr_clock_bridge_m1_writedata /= tse_ddr_clock_bridge_m1_writedata_last_time)))) AND tse_ddr_clock_bridge_m1_write)) = '1' then 
          write(write_line62, now);
          write(write_line62, string'(": "));
          write(write_line62, string'("tse_ddr_clock_bridge_m1_writedata did not heed wait!!!"));
          write(output, write_line62.all);
          deallocate (write_line62);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo read when empty, which is an e_process
    process (clk)
    VARIABLE write_line63 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((empty_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo AND read_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo)) = '1' then 
          write(write_line63, now);
          write(write_line63, string'(": "));
          write(write_line63, string'("tse_ddr_clock_bridge/m1 negative rdv fifo selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo: read AND empty."));
          write(output, write_line63.all & CR);
          deallocate (write_line63);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo write when full, which is an e_process
    process (clk)
    VARIABLE write_line64 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((full_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo AND write_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo) AND NOT read_selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo)) = '1' then 
          write(write_line64, now);
          write(write_line64, string'(": "));
          write(write_line64, string'("tse_ddr_clock_bridge/m1 negative rdv fifo selecto_nrdv_tse_ddr_clock_bridge_m1_1_sdram_s1_fifo: write AND full."));
          write(output, write_line64.all & CR);
          deallocate (write_line64);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tse_ddr_clock_bridge_bridge_arbitrator is 
end entity tse_ddr_clock_bridge_bridge_arbitrator;


architecture europa of tse_ddr_clock_bridge_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tse_mac_control_port_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                 signal cpuNios_data_master_read : IN STD_LOGIC;
                 signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                 signal cpuNios_data_master_write : IN STD_LOGIC;
                 signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal tse_mac_control_port_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_control_port_waitrequest : IN STD_LOGIC;

              -- outputs:
                 signal cpuNios_data_master_granted_tse_mac_control_port : OUT STD_LOGIC;
                 signal cpuNios_data_master_qualified_request_tse_mac_control_port : OUT STD_LOGIC;
                 signal cpuNios_data_master_read_data_valid_tse_mac_control_port : OUT STD_LOGIC;
                 signal cpuNios_data_master_requests_tse_mac_control_port : OUT STD_LOGIC;
                 signal d1_tse_mac_control_port_end_xfer : OUT STD_LOGIC;
                 signal tse_mac_control_port_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal tse_mac_control_port_read : OUT STD_LOGIC;
                 signal tse_mac_control_port_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_control_port_reset : OUT STD_LOGIC;
                 signal tse_mac_control_port_waitrequest_from_sa : OUT STD_LOGIC;
                 signal tse_mac_control_port_write : OUT STD_LOGIC;
                 signal tse_mac_control_port_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity tse_mac_control_port_arbitrator;


architecture europa of tse_mac_control_port_arbitrator is
                signal cpuNios_data_master_arbiterlock :  STD_LOGIC;
                signal cpuNios_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpuNios_data_master_continuerequest :  STD_LOGIC;
                signal cpuNios_data_master_saved_grant_tse_mac_control_port :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_tse_mac_control_port :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpuNios_data_master_granted_tse_mac_control_port :  STD_LOGIC;
                signal internal_cpuNios_data_master_qualified_request_tse_mac_control_port :  STD_LOGIC;
                signal internal_cpuNios_data_master_requests_tse_mac_control_port :  STD_LOGIC;
                signal internal_tse_mac_control_port_waitrequest_from_sa :  STD_LOGIC;
                signal shifted_address_to_tse_mac_control_port_from_cpuNios_data_master :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal tse_mac_control_port_allgrants :  STD_LOGIC;
                signal tse_mac_control_port_allow_new_arb_cycle :  STD_LOGIC;
                signal tse_mac_control_port_any_bursting_master_saved_grant :  STD_LOGIC;
                signal tse_mac_control_port_any_continuerequest :  STD_LOGIC;
                signal tse_mac_control_port_arb_counter_enable :  STD_LOGIC;
                signal tse_mac_control_port_arb_share_counter :  STD_LOGIC;
                signal tse_mac_control_port_arb_share_counter_next_value :  STD_LOGIC;
                signal tse_mac_control_port_arb_share_set_values :  STD_LOGIC;
                signal tse_mac_control_port_beginbursttransfer_internal :  STD_LOGIC;
                signal tse_mac_control_port_begins_xfer :  STD_LOGIC;
                signal tse_mac_control_port_end_xfer :  STD_LOGIC;
                signal tse_mac_control_port_firsttransfer :  STD_LOGIC;
                signal tse_mac_control_port_grant_vector :  STD_LOGIC;
                signal tse_mac_control_port_in_a_read_cycle :  STD_LOGIC;
                signal tse_mac_control_port_in_a_write_cycle :  STD_LOGIC;
                signal tse_mac_control_port_master_qreq_vector :  STD_LOGIC;
                signal tse_mac_control_port_non_bursting_master_requests :  STD_LOGIC;
                signal tse_mac_control_port_reg_firsttransfer :  STD_LOGIC;
                signal tse_mac_control_port_slavearbiterlockenable :  STD_LOGIC;
                signal tse_mac_control_port_slavearbiterlockenable2 :  STD_LOGIC;
                signal tse_mac_control_port_unreg_firsttransfer :  STD_LOGIC;
                signal tse_mac_control_port_waits_for_read :  STD_LOGIC;
                signal tse_mac_control_port_waits_for_write :  STD_LOGIC;
                signal wait_for_tse_mac_control_port_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT tse_mac_control_port_end_xfer;
    end if;

  end process;

  tse_mac_control_port_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpuNios_data_master_qualified_request_tse_mac_control_port);
  --assign tse_mac_control_port_readdata_from_sa = tse_mac_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  tse_mac_control_port_readdata_from_sa <= tse_mac_control_port_readdata;
  internal_cpuNios_data_master_requests_tse_mac_control_port <= to_std_logic(((Std_Logic_Vector'(cpuNios_data_master_address_to_slave(26 DOWNTO 10) & std_logic_vector'("0000000000")) = std_logic_vector'("100000000000100000000000000")))) AND ((cpuNios_data_master_read OR cpuNios_data_master_write));
  --assign tse_mac_control_port_waitrequest_from_sa = tse_mac_control_port_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_tse_mac_control_port_waitrequest_from_sa <= tse_mac_control_port_waitrequest;
  --tse_mac_control_port_arb_share_counter set values, which is an e_mux
  tse_mac_control_port_arb_share_set_values <= std_logic'('1');
  --tse_mac_control_port_non_bursting_master_requests mux, which is an e_mux
  tse_mac_control_port_non_bursting_master_requests <= internal_cpuNios_data_master_requests_tse_mac_control_port;
  --tse_mac_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  tse_mac_control_port_any_bursting_master_saved_grant <= std_logic'('0');
  --tse_mac_control_port_arb_share_counter_next_value assignment, which is an e_assign
  tse_mac_control_port_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(tse_mac_control_port_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_mac_control_port_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(tse_mac_control_port_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_mac_control_port_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --tse_mac_control_port_allgrants all slave grants, which is an e_mux
  tse_mac_control_port_allgrants <= tse_mac_control_port_grant_vector;
  --tse_mac_control_port_end_xfer assignment, which is an e_assign
  tse_mac_control_port_end_xfer <= NOT ((tse_mac_control_port_waits_for_read OR tse_mac_control_port_waits_for_write));
  --end_xfer_arb_share_counter_term_tse_mac_control_port arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_tse_mac_control_port <= tse_mac_control_port_end_xfer AND (((NOT tse_mac_control_port_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --tse_mac_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  tse_mac_control_port_arb_counter_enable <= ((end_xfer_arb_share_counter_term_tse_mac_control_port AND tse_mac_control_port_allgrants)) OR ((end_xfer_arb_share_counter_term_tse_mac_control_port AND NOT tse_mac_control_port_non_bursting_master_requests));
  --tse_mac_control_port_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_mac_control_port_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(tse_mac_control_port_arb_counter_enable) = '1' then 
        tse_mac_control_port_arb_share_counter <= tse_mac_control_port_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --tse_mac_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_mac_control_port_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((tse_mac_control_port_master_qreq_vector AND end_xfer_arb_share_counter_term_tse_mac_control_port)) OR ((end_xfer_arb_share_counter_term_tse_mac_control_port AND NOT tse_mac_control_port_non_bursting_master_requests)))) = '1' then 
        tse_mac_control_port_slavearbiterlockenable <= tse_mac_control_port_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpuNios/data_master tse_mac/control_port arbiterlock, which is an e_assign
  cpuNios_data_master_arbiterlock <= tse_mac_control_port_slavearbiterlockenable AND cpuNios_data_master_continuerequest;
  --tse_mac_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  tse_mac_control_port_slavearbiterlockenable2 <= tse_mac_control_port_arb_share_counter_next_value;
  --cpuNios/data_master tse_mac/control_port arbiterlock2, which is an e_assign
  cpuNios_data_master_arbiterlock2 <= tse_mac_control_port_slavearbiterlockenable2 AND cpuNios_data_master_continuerequest;
  --tse_mac_control_port_any_continuerequest at least one master continues requesting, which is an e_assign
  tse_mac_control_port_any_continuerequest <= std_logic'('1');
  --cpuNios_data_master_continuerequest continued request, which is an e_assign
  cpuNios_data_master_continuerequest <= std_logic'('1');
  internal_cpuNios_data_master_qualified_request_tse_mac_control_port <= internal_cpuNios_data_master_requests_tse_mac_control_port AND NOT ((((cpuNios_data_master_read AND (NOT cpuNios_data_master_waitrequest))) OR (((NOT cpuNios_data_master_waitrequest) AND cpuNios_data_master_write))));
  --tse_mac_control_port_writedata mux, which is an e_mux
  tse_mac_control_port_writedata <= cpuNios_data_master_writedata;
  --master is always granted when requested
  internal_cpuNios_data_master_granted_tse_mac_control_port <= internal_cpuNios_data_master_qualified_request_tse_mac_control_port;
  --cpuNios/data_master saved-grant tse_mac/control_port, which is an e_assign
  cpuNios_data_master_saved_grant_tse_mac_control_port <= internal_cpuNios_data_master_requests_tse_mac_control_port;
  --allow new arb cycle for tse_mac/control_port, which is an e_assign
  tse_mac_control_port_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  tse_mac_control_port_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  tse_mac_control_port_master_qreq_vector <= std_logic'('1');
  --~tse_mac_control_port_reset assignment, which is an e_assign
  tse_mac_control_port_reset <= NOT reset_n;
  --tse_mac_control_port_firsttransfer first transaction, which is an e_assign
  tse_mac_control_port_firsttransfer <= A_WE_StdLogic((std_logic'(tse_mac_control_port_begins_xfer) = '1'), tse_mac_control_port_unreg_firsttransfer, tse_mac_control_port_reg_firsttransfer);
  --tse_mac_control_port_unreg_firsttransfer first transaction, which is an e_assign
  tse_mac_control_port_unreg_firsttransfer <= NOT ((tse_mac_control_port_slavearbiterlockenable AND tse_mac_control_port_any_continuerequest));
  --tse_mac_control_port_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_mac_control_port_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(tse_mac_control_port_begins_xfer) = '1' then 
        tse_mac_control_port_reg_firsttransfer <= tse_mac_control_port_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --tse_mac_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  tse_mac_control_port_beginbursttransfer_internal <= tse_mac_control_port_begins_xfer;
  --tse_mac_control_port_read assignment, which is an e_mux
  tse_mac_control_port_read <= internal_cpuNios_data_master_granted_tse_mac_control_port AND cpuNios_data_master_read;
  --tse_mac_control_port_write assignment, which is an e_mux
  tse_mac_control_port_write <= internal_cpuNios_data_master_granted_tse_mac_control_port AND cpuNios_data_master_write;
  shifted_address_to_tse_mac_control_port_from_cpuNios_data_master <= cpuNios_data_master_address_to_slave;
  --tse_mac_control_port_address mux, which is an e_mux
  tse_mac_control_port_address <= A_EXT (A_SRL(shifted_address_to_tse_mac_control_port_from_cpuNios_data_master,std_logic_vector'("00000000000000000000000000000010")), 8);
  --d1_tse_mac_control_port_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_tse_mac_control_port_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_tse_mac_control_port_end_xfer <= tse_mac_control_port_end_xfer;
    end if;

  end process;

  --tse_mac_control_port_waits_for_read in a cycle, which is an e_mux
  tse_mac_control_port_waits_for_read <= tse_mac_control_port_in_a_read_cycle AND internal_tse_mac_control_port_waitrequest_from_sa;
  --tse_mac_control_port_in_a_read_cycle assignment, which is an e_assign
  tse_mac_control_port_in_a_read_cycle <= internal_cpuNios_data_master_granted_tse_mac_control_port AND cpuNios_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= tse_mac_control_port_in_a_read_cycle;
  --tse_mac_control_port_waits_for_write in a cycle, which is an e_mux
  tse_mac_control_port_waits_for_write <= tse_mac_control_port_in_a_write_cycle AND internal_tse_mac_control_port_waitrequest_from_sa;
  --tse_mac_control_port_in_a_write_cycle assignment, which is an e_assign
  tse_mac_control_port_in_a_write_cycle <= internal_cpuNios_data_master_granted_tse_mac_control_port AND cpuNios_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= tse_mac_control_port_in_a_write_cycle;
  wait_for_tse_mac_control_port_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpuNios_data_master_granted_tse_mac_control_port <= internal_cpuNios_data_master_granted_tse_mac_control_port;
  --vhdl renameroo for output signals
  cpuNios_data_master_qualified_request_tse_mac_control_port <= internal_cpuNios_data_master_qualified_request_tse_mac_control_port;
  --vhdl renameroo for output signals
  cpuNios_data_master_requests_tse_mac_control_port <= internal_cpuNios_data_master_requests_tse_mac_control_port;
  --vhdl renameroo for output signals
  tse_mac_control_port_waitrequest_from_sa <= internal_tse_mac_control_port_waitrequest_from_sa;
--synthesis translate_off
    --tse_mac/control_port enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tse_mac_transmit_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sgdma_tx_out_endofpacket : IN STD_LOGIC;
                 signal sgdma_tx_out_error : IN STD_LOGIC;
                 signal sgdma_tx_out_startofpacket : IN STD_LOGIC;
                 signal sgdma_tx_out_valid : IN STD_LOGIC;
                 signal tse_mac_transmit_ready : IN STD_LOGIC;

              -- outputs:
                 signal tse_mac_transmit_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_transmit_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal tse_mac_transmit_endofpacket : OUT STD_LOGIC;
                 signal tse_mac_transmit_error : OUT STD_LOGIC;
                 signal tse_mac_transmit_ready_from_sa : OUT STD_LOGIC;
                 signal tse_mac_transmit_startofpacket : OUT STD_LOGIC;
                 signal tse_mac_transmit_valid : OUT STD_LOGIC
              );
end entity tse_mac_transmit_arbitrator;


architecture europa of tse_mac_transmit_arbitrator is

begin

  --mux tse_mac_transmit_data, which is an e_mux
  tse_mac_transmit_data <= sgdma_tx_out_data;
  --mux tse_mac_transmit_endofpacket, which is an e_mux
  tse_mac_transmit_endofpacket <= sgdma_tx_out_endofpacket;
  --mux tse_mac_transmit_error, which is an e_mux
  tse_mac_transmit_error <= sgdma_tx_out_error;
  --mux tse_mac_transmit_empty, which is an e_mux
  tse_mac_transmit_empty <= sgdma_tx_out_empty;
  --assign tse_mac_transmit_ready_from_sa = tse_mac_transmit_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  tse_mac_transmit_ready_from_sa <= tse_mac_transmit_ready;
  --mux tse_mac_transmit_startofpacket, which is an e_mux
  tse_mac_transmit_startofpacket <= sgdma_tx_out_startofpacket;
  --mux tse_mac_transmit_valid, which is an e_mux
  tse_mac_transmit_valid <= sgdma_tx_out_valid;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tse_mac_receive_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_in_ready_from_sa : IN STD_LOGIC;
                 signal tse_mac_receive_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_receive_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal tse_mac_receive_endofpacket : IN STD_LOGIC;
                 signal tse_mac_receive_error : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal tse_mac_receive_startofpacket : IN STD_LOGIC;
                 signal tse_mac_receive_valid : IN STD_LOGIC;

              -- outputs:
                 signal tse_mac_receive_ready : OUT STD_LOGIC
              );
end entity tse_mac_receive_arbitrator;


architecture europa of tse_mac_receive_arbitrator is

begin

  --mux tse_mac_receive_ready, which is an e_mux
  tse_mac_receive_ready <= sgdma_rx_in_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity processador_reset_clk100MHz_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity processador_reset_clk100MHz_domain_synch_module;


architecture europa of processador_reset_clk100MHz_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity processador_reset_sdram_phy_clk_out_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity processador_reset_sdram_phy_clk_out_domain_synch_module;


architecture europa of processador_reset_sdram_phy_clk_out_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity processador is 
        port (
              -- 1) global signals:
                 signal clk100MHz : IN STD_LOGIC;
                 signal clk50Mhz : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_aux_full_rate_clk_out : OUT STD_LOGIC;
                 signal sdram_aux_half_rate_clk_out : OUT STD_LOGIC;
                 signal sdram_phy_clk_out : OUT STD_LOGIC;

              -- the_fft_pipeline_0
                 signal counter_from_the_fft_pipeline_0 : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                 signal rx_in_to_the_fft_pipeline_0 : IN STD_LOGIC;
                 signal tx_out_from_the_fft_pipeline_0 : OUT STD_LOGIC;

              -- the_lcd_i2c_en
                 signal out_port_from_the_lcd_i2c_en : OUT STD_LOGIC;

              -- the_lcd_i2c_scl
                 signal out_port_from_the_lcd_i2c_scl : OUT STD_LOGIC;

              -- the_lcd_i2c_sdat
                 signal bidir_port_to_and_from_the_lcd_i2c_sdat : INOUT STD_LOGIC;

              -- the_lcd_sync_generator
                 signal DEN_from_the_lcd_sync_generator : OUT STD_LOGIC;
                 signal HD_from_the_lcd_sync_generator : OUT STD_LOGIC;
                 signal RGB_OUT_from_the_lcd_sync_generator : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal VD_from_the_lcd_sync_generator : OUT STD_LOGIC;

              -- the_sdram
                 signal global_reset_n_to_the_sdram : IN STD_LOGIC;
                 signal local_init_done_from_the_sdram : OUT STD_LOGIC;
                 signal local_refresh_ack_from_the_sdram : OUT STD_LOGIC;
                 signal local_wdata_req_from_the_sdram : OUT STD_LOGIC;
                 signal mem_addr_from_the_sdram : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal mem_ba_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal mem_cas_n_from_the_sdram : OUT STD_LOGIC;
                 signal mem_cke_from_the_sdram : OUT STD_LOGIC;
                 signal mem_clk_n_to_and_from_the_sdram : INOUT STD_LOGIC;
                 signal mem_clk_to_and_from_the_sdram : INOUT STD_LOGIC;
                 signal mem_cs_n_from_the_sdram : OUT STD_LOGIC;
                 signal mem_dm_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal mem_dq_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal mem_dqs_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal mem_ras_n_from_the_sdram : OUT STD_LOGIC;
                 signal mem_we_n_from_the_sdram : OUT STD_LOGIC;
                 signal reset_phy_clk_n_from_the_sdram : OUT STD_LOGIC;

              -- the_tse_mac
                 signal ena_10_from_the_tse_mac : OUT STD_LOGIC;
                 signal eth_mode_from_the_tse_mac : OUT STD_LOGIC;
                 signal gm_rx_d_to_the_tse_mac : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gm_rx_dv_to_the_tse_mac : IN STD_LOGIC;
                 signal gm_rx_err_to_the_tse_mac : IN STD_LOGIC;
                 signal gm_tx_d_from_the_tse_mac : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gm_tx_en_from_the_tse_mac : OUT STD_LOGIC;
                 signal gm_tx_err_from_the_tse_mac : OUT STD_LOGIC;
                 signal m_rx_col_to_the_tse_mac : IN STD_LOGIC;
                 signal m_rx_crs_to_the_tse_mac : IN STD_LOGIC;
                 signal m_rx_d_to_the_tse_mac : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal m_rx_en_to_the_tse_mac : IN STD_LOGIC;
                 signal m_rx_err_to_the_tse_mac : IN STD_LOGIC;
                 signal m_tx_d_from_the_tse_mac : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal m_tx_en_from_the_tse_mac : OUT STD_LOGIC;
                 signal m_tx_err_from_the_tse_mac : OUT STD_LOGIC;
                 signal mdc_from_the_tse_mac : OUT STD_LOGIC;
                 signal mdio_in_to_the_tse_mac : IN STD_LOGIC;
                 signal mdio_oen_from_the_tse_mac : OUT STD_LOGIC;
                 signal mdio_out_from_the_tse_mac : OUT STD_LOGIC;
                 signal rx_clk_to_the_tse_mac : IN STD_LOGIC;
                 signal set_1000_to_the_tse_mac : IN STD_LOGIC;
                 signal set_10_to_the_tse_mac : IN STD_LOGIC;
                 signal tx_clk_to_the_tse_mac : IN STD_LOGIC
              );
end entity processador;


architecture europa of processador is
component cpuNios_jtag_debug_module_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpuNios_data_master_debugaccess : IN STD_LOGIC;
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpuNios_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_instruction_master_read : IN STD_LOGIC;
                    signal cpuNios_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpuNios_jtag_debug_module_resetrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_granted_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                    signal cpuNios_instruction_master_granted_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                    signal cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                    signal cpuNios_instruction_master_read_data_valid_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                    signal cpuNios_instruction_master_requests_cpuNios_jtag_debug_module : OUT STD_LOGIC;
                    signal cpuNios_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal cpuNios_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                    signal cpuNios_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpuNios_jtag_debug_module_chipselect : OUT STD_LOGIC;
                    signal cpuNios_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                    signal cpuNios_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpuNios_jtag_debug_module_reset_n : OUT STD_LOGIC;
                    signal cpuNios_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                    signal cpuNios_jtag_debug_module_write : OUT STD_LOGIC;
                    signal cpuNios_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpuNios_jtag_debug_module_end_xfer : OUT STD_LOGIC
                 );
end component cpuNios_jtag_debug_module_arbitrator;

component cpuNios_data_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clk100MHz : IN STD_LOGIC;
                    signal clk100MHz_reset_n : IN STD_LOGIC;
                    signal cpuNios_data_master_address : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_granted_cpuNios_jtag_debug_module : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_descriptor_memory_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_lcd_i2c_en_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_lcd_i2c_scl_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_lcd_i2c_sdat_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_performance_counter_control_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_sgdma_rx_csr : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_sgdma_tx_csr : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_sysid_control_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_granted_tse_mac_control_port : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_lcd_i2c_en_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_performance_counter_control_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_sgdma_rx_csr : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_sgdma_tx_csr : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_sysid_control_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_tse_mac_control_port : IN STD_LOGIC;
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_cpuNios_jtag_debug_module : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_fft_pipeline_0_avalon_slave_0 : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_lcd_i2c_en_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_lcd_i2c_scl_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_lcd_i2c_sdat_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_performance_counter_control_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_sgdma_rx_csr : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_sgdma_tx_csr : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_tse_mac_control_port : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_cpuNios_jtag_debug_module : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_descriptor_memory_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_lcd_i2c_en_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_lcd_i2c_scl_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_lcd_i2c_sdat_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_performance_counter_control_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_sgdma_rx_csr : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_sgdma_tx_csr : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_sysid_control_slave : IN STD_LOGIC;
                    signal cpuNios_data_master_requests_tse_mac_control_port : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal d1_cpuNios_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_cpu_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                    signal d1_fft_pipeline_0_avalon_slave_0_end_xfer : IN STD_LOGIC;
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                    signal d1_lcd_i2c_en_s1_end_xfer : IN STD_LOGIC;
                    signal d1_lcd_i2c_scl_s1_end_xfer : IN STD_LOGIC;
                    signal d1_lcd_i2c_sdat_s1_end_xfer : IN STD_LOGIC;
                    signal d1_performance_counter_control_slave_end_xfer : IN STD_LOGIC;
                    signal d1_sgdma_rx_csr_end_xfer : IN STD_LOGIC;
                    signal d1_sgdma_tx_csr_end_xfer : IN STD_LOGIC;
                    signal d1_sys_clk_timer_s1_end_xfer : IN STD_LOGIC;
                    signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                    signal d1_tse_mac_control_port_end_xfer : IN STD_LOGIC;
                    signal descriptor_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal fft_pipeline_0_avalon_slave_0_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal lcd_i2c_en_s1_readdata_from_sa : IN STD_LOGIC;
                    signal lcd_i2c_scl_s1_readdata_from_sa : IN STD_LOGIC;
                    signal lcd_i2c_sdat_s1_readdata_from_sa : IN STD_LOGIC;
                    signal lcd_sgdma_csr_irq_from_sa : IN STD_LOGIC;
                    signal performance_counter_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                    signal registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_csr_irq_from_sa : IN STD_LOGIC;
                    signal sgdma_rx_csr_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_csr_irq_from_sa : IN STD_LOGIC;
                    signal sgdma_tx_csr_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sys_clk_timer_s1_irq_from_sa : IN STD_LOGIC;
                    signal sys_clk_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_control_port_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpuNios_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpuNios_data_master_waitrequest : OUT STD_LOGIC
                 );
end component cpuNios_data_master_arbitrator;

component cpuNios_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_instruction_master_address : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_instruction_master_granted_cpuNios_jtag_debug_module : IN STD_LOGIC;
                    signal cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module : IN STD_LOGIC;
                    signal cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpuNios_instruction_master_read : IN STD_LOGIC;
                    signal cpuNios_instruction_master_read_data_valid_cpuNios_jtag_debug_module : IN STD_LOGIC;
                    signal cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpuNios_instruction_master_requests_cpuNios_jtag_debug_module : IN STD_LOGIC;
                    signal cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal cpuNios_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal d1_cpuNios_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_cpu_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpuNios_instruction_master_waitrequest : OUT STD_LOGIC
                 );
end component cpuNios_instruction_master_arbitrator;

component cpuNios is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d_irq : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_waitrequest : IN STD_LOGIC;
                    signal i_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_waitrequest : IN STD_LOGIC;
                    signal jtag_debug_module_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal jtag_debug_module_begintransfer : IN STD_LOGIC;
                    signal jtag_debug_module_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal jtag_debug_module_debugaccess : IN STD_LOGIC;
                    signal jtag_debug_module_select : IN STD_LOGIC;
                    signal jtag_debug_module_write : IN STD_LOGIC;
                    signal jtag_debug_module_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d_address : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal d_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_read : OUT STD_LOGIC;
                    signal d_write : OUT STD_LOGIC;
                    signal d_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_address : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal i_read : OUT STD_LOGIC;
                    signal jtag_debug_module_debugaccess_to_roms : OUT STD_LOGIC;
                    signal jtag_debug_module_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_debug_module_resetrequest : OUT STD_LOGIC
                 );
end component cpuNios;

component cpu_ddr_clock_bridge_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpuNios_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_instruction_master_read : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_endofpacket : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_readdatavalid : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_read : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_s1_reset_n : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_write : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_ddr_clock_bridge_s1_end_xfer : OUT STD_LOGIC
                 );
end component cpu_ddr_clock_bridge_s1_arbitrator;

component cpu_ddr_clock_bridge_m1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_granted_sdram_s1 : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_requests_sdram_s1 : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_lcd_sgdma_csr_end_xfer : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal lcd_sgdma_csr_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_ddr_clock_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_latency_counter : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_readdatavalid : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_reset_n : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_waitrequest : OUT STD_LOGIC
                 );
end component cpu_ddr_clock_bridge_m1_arbitrator;

component cpu_ddr_clock_bridge is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_readdatavalid : IN STD_LOGIC;
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_readdatavalid : OUT STD_LOGIC;
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component cpu_ddr_clock_bridge;

component cpu_ddr_clock_bridge_bridge_arbitrator is 
end component cpu_ddr_clock_bridge_bridge_arbitrator;

component descriptor_memory_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_burstcount : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_chipselect : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_dbs_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_dbs_write_32 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_read : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal d1_descriptor_memory_s1_end_xfer : OUT STD_LOGIC;
                    signal descriptor_memory_s1_address : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal descriptor_memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal descriptor_memory_s1_chipselect : OUT STD_LOGIC;
                    signal descriptor_memory_s1_clken : OUT STD_LOGIC;
                    signal descriptor_memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_memory_s1_reset : OUT STD_LOGIC;
                    signal descriptor_memory_s1_write : OUT STD_LOGIC;
                    signal descriptor_memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1 : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_m1_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC
                 );
end component descriptor_memory_s1_arbitrator;

component descriptor_memory is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clken : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component descriptor_memory;

component descriptor_offset_bridge_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal descriptor_offset_bridge_s1_endofpacket : IN STD_LOGIC;
                    signal descriptor_offset_bridge_s1_readdata : IN STD_LOGIC_VECTOR (255 DOWNTO 0);
                    signal descriptor_offset_bridge_s1_readdatavalid : IN STD_LOGIC;
                    signal descriptor_offset_bridge_s1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_read_latency_counter : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_read : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_write_write : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_read_latency_counter : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_read : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_write_write : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal d1_descriptor_offset_bridge_s1_end_xfer : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal descriptor_offset_bridge_s1_arbiterlock : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_arbiterlock2 : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_burstcount : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_offset_bridge_s1_chipselect : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_debugaccess : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal descriptor_offset_bridge_s1_read : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (255 DOWNTO 0);
                    signal descriptor_offset_bridge_s1_reset_n : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_write : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (255 DOWNTO 0);
                    signal sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 : OUT STD_LOGIC
                 );
end component descriptor_offset_bridge_s1_arbitrator;

component descriptor_offset_bridge_m1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                    signal descriptor_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_address : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_burstcount : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1 : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_chipselect : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_granted_descriptor_memory_s1 : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_read : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_requests_descriptor_memory_s1 : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_write : IN STD_LOGIC;
                    signal descriptor_offset_bridge_m1_writedata : IN STD_LOGIC_VECTOR (255 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal descriptor_offset_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_dbs_address : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_dbs_write_32 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_latency_counter : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (255 DOWNTO 0);
                    signal descriptor_offset_bridge_m1_readdatavalid : OUT STD_LOGIC;
                    signal descriptor_offset_bridge_m1_waitrequest : OUT STD_LOGIC
                 );
end component descriptor_offset_bridge_m1_arbitrator;

component descriptor_offset_bridge is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal m1_endofpacket : IN STD_LOGIC;
                    signal m1_readdata : IN STD_LOGIC_VECTOR (255 DOWNTO 0);
                    signal m1_readdatavalid : IN STD_LOGIC;
                    signal m1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal s1_address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal s1_arbiterlock : IN STD_LOGIC;
                    signal s1_arbiterlock2 : IN STD_LOGIC;
                    signal s1_burstcount : IN STD_LOGIC;
                    signal s1_byteenable : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal s1_chipselect : IN STD_LOGIC;
                    signal s1_debugaccess : IN STD_LOGIC;
                    signal s1_nativeaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal s1_read : IN STD_LOGIC;
                    signal s1_write : IN STD_LOGIC;
                    signal s1_writedata : IN STD_LOGIC_VECTOR (255 DOWNTO 0);

                 -- outputs:
                    signal m1_address : OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal m1_burstcount : OUT STD_LOGIC;
                    signal m1_byteenable : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m1_chipselect : OUT STD_LOGIC;
                    signal m1_debugaccess : OUT STD_LOGIC;
                    signal m1_read : OUT STD_LOGIC;
                    signal m1_write : OUT STD_LOGIC;
                    signal m1_writedata : OUT STD_LOGIC_VECTOR (255 DOWNTO 0);
                    signal s1_endofpacket : OUT STD_LOGIC;
                    signal s1_readdata : OUT STD_LOGIC_VECTOR (255 DOWNTO 0);
                    signal s1_readdatavalid : OUT STD_LOGIC;
                    signal s1_waitrequest : OUT STD_LOGIC
                 );
end component descriptor_offset_bridge;

component descriptor_offset_bridge_bridge_arbitrator is 
end component descriptor_offset_bridge_bridge_arbitrator;

component fft_pipeline_0_avalon_slave_0_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal fft_pipeline_0_avalon_slave_0_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_fft_pipeline_0_avalon_slave_0 : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 : OUT STD_LOGIC;
                    signal d1_fft_pipeline_0_avalon_slave_0_end_xfer : OUT STD_LOGIC;
                    signal fft_pipeline_0_avalon_slave_0_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal fft_pipeline_0_avalon_slave_0_chipselect : OUT STD_LOGIC;
                    signal fft_pipeline_0_avalon_slave_0_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal fft_pipeline_0_avalon_slave_0_reset : OUT STD_LOGIC;
                    signal fft_pipeline_0_avalon_slave_0_write : OUT STD_LOGIC;
                    signal fft_pipeline_0_avalon_slave_0_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component fft_pipeline_0_avalon_slave_0_arbitrator;

component fft_pipeline_0 is 
           port (
                 -- inputs:
                    signal addr : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal clr_n : IN STD_LOGIC;
                    signal cs : IN STD_LOGIC;
                    signal rx_in : IN STD_LOGIC;
                    signal wr : IN STD_LOGIC;
                    signal wr_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal counter : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal rd_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tx_out : OUT STD_LOGIC
                 );
end component fft_pipeline_0;

component jtag_uart_avalon_jtag_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component jtag_uart_avalon_jtag_slave_arbitrator;

component jtag_uart is 
           port (
                 -- inputs:
                    signal av_address : IN STD_LOGIC;
                    signal av_chipselect : IN STD_LOGIC;
                    signal av_read_n : IN STD_LOGIC;
                    signal av_write_n : IN STD_LOGIC;
                    signal av_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_irq : OUT STD_LOGIC;
                    signal av_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_waitrequest : OUT STD_LOGIC;
                    signal dataavailable : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component jtag_uart;

component lcd_24_to_8_bits_dfa_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_in_ready : IN STD_LOGIC;
                    signal lcd_pixel_converter_out_data : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal lcd_pixel_converter_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_pixel_converter_out_endofpacket : IN STD_LOGIC;
                    signal lcd_pixel_converter_out_startofpacket : IN STD_LOGIC;
                    signal lcd_pixel_converter_out_valid : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_24_to_8_bits_dfa_in_data : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal lcd_24_to_8_bits_dfa_in_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_24_to_8_bits_dfa_in_endofpacket : OUT STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_in_ready_from_sa : OUT STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_in_reset_n : OUT STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_in_startofpacket : OUT STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_in_valid : OUT STD_LOGIC
                 );
end component lcd_24_to_8_bits_dfa_in_arbitrator;

component lcd_24_to_8_bits_dfa_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_out_data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal lcd_24_to_8_bits_dfa_out_empty : IN STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_out_endofpacket : IN STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_out_startofpacket : IN STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_out_valid : IN STD_LOGIC;
                    signal lcd_sync_generator_in_ready_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_24_to_8_bits_dfa_out_ready : OUT STD_LOGIC
                 );
end component lcd_24_to_8_bits_dfa_out_arbitrator;

component lcd_24_to_8_bits_dfa is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal in_data : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal in_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal in_endofpacket : IN STD_LOGIC;
                    signal in_startofpacket : IN STD_LOGIC;
                    signal in_valid : IN STD_LOGIC;
                    signal out_ready : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal in_ready : OUT STD_LOGIC;
                    signal out_data : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal out_empty : OUT STD_LOGIC;
                    signal out_endofpacket : OUT STD_LOGIC;
                    signal out_startofpacket : OUT STD_LOGIC;
                    signal out_valid : OUT STD_LOGIC
                 );
end component lcd_24_to_8_bits_dfa;

component lcd_64_to_32_bits_dfa_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_in_ready : IN STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_ta_fifo_to_dfa_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_ta_fifo_to_dfa_out_endofpacket : IN STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_out_startofpacket : IN STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_out_valid : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_64_to_32_bits_dfa_in_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_64_to_32_bits_dfa_in_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_64_to_32_bits_dfa_in_endofpacket : OUT STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_in_ready_from_sa : OUT STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_in_reset_n : OUT STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_in_startofpacket : OUT STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_in_valid : OUT STD_LOGIC
                 );
end component lcd_64_to_32_bits_dfa_in_arbitrator;

component lcd_64_to_32_bits_dfa_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_64_to_32_bits_dfa_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_64_to_32_bits_dfa_out_endofpacket : IN STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_out_startofpacket : IN STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_out_valid : IN STD_LOGIC;
                    signal lcd_pixel_converter_in_ready_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_64_to_32_bits_dfa_out_ready : OUT STD_LOGIC
                 );
end component lcd_64_to_32_bits_dfa_out_arbitrator;

component lcd_64_to_32_bits_dfa is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal in_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal in_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal in_endofpacket : IN STD_LOGIC;
                    signal in_startofpacket : IN STD_LOGIC;
                    signal in_valid : IN STD_LOGIC;
                    signal out_ready : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal in_ready : OUT STD_LOGIC;
                    signal out_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal out_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal out_endofpacket : OUT STD_LOGIC;
                    signal out_startofpacket : OUT STD_LOGIC;
                    signal out_valid : OUT STD_LOGIC
                 );
end component lcd_64_to_32_bits_dfa;

component lcd_i2c_en_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_i2c_en_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_granted_lcd_i2c_en_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_lcd_i2c_en_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_lcd_i2c_en_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_lcd_i2c_en_s1 : OUT STD_LOGIC;
                    signal d1_lcd_i2c_en_s1_end_xfer : OUT STD_LOGIC;
                    signal lcd_i2c_en_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_i2c_en_s1_chipselect : OUT STD_LOGIC;
                    signal lcd_i2c_en_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal lcd_i2c_en_s1_reset_n : OUT STD_LOGIC;
                    signal lcd_i2c_en_s1_write_n : OUT STD_LOGIC;
                    signal lcd_i2c_en_s1_writedata : OUT STD_LOGIC
                 );
end component lcd_i2c_en_s1_arbitrator;

component lcd_i2c_en is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component lcd_i2c_en;

component lcd_i2c_scl_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_i2c_scl_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_granted_lcd_i2c_scl_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_lcd_i2c_scl_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_lcd_i2c_scl_s1 : OUT STD_LOGIC;
                    signal d1_lcd_i2c_scl_s1_end_xfer : OUT STD_LOGIC;
                    signal lcd_i2c_scl_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_i2c_scl_s1_chipselect : OUT STD_LOGIC;
                    signal lcd_i2c_scl_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal lcd_i2c_scl_s1_reset_n : OUT STD_LOGIC;
                    signal lcd_i2c_scl_s1_write_n : OUT STD_LOGIC;
                    signal lcd_i2c_scl_s1_writedata : OUT STD_LOGIC
                 );
end component lcd_i2c_scl_s1_arbitrator;

component lcd_i2c_scl is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component lcd_i2c_scl;

component lcd_i2c_sdat_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_i2c_sdat_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_granted_lcd_i2c_sdat_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_lcd_i2c_sdat_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_lcd_i2c_sdat_s1 : OUT STD_LOGIC;
                    signal d1_lcd_i2c_sdat_s1_end_xfer : OUT STD_LOGIC;
                    signal lcd_i2c_sdat_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_i2c_sdat_s1_chipselect : OUT STD_LOGIC;
                    signal lcd_i2c_sdat_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal lcd_i2c_sdat_s1_reset_n : OUT STD_LOGIC;
                    signal lcd_i2c_sdat_s1_write_n : OUT STD_LOGIC;
                    signal lcd_i2c_sdat_s1_writedata : OUT STD_LOGIC
                 );
end component lcd_i2c_sdat_s1_arbitrator;

component lcd_i2c_sdat is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal bidir_port : INOUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component lcd_i2c_sdat;

component lcd_pixel_converter_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_64_to_32_bits_dfa_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_64_to_32_bits_dfa_out_endofpacket : IN STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_out_startofpacket : IN STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_out_valid : IN STD_LOGIC;
                    signal lcd_pixel_converter_in_ready : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_pixel_converter_in_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_pixel_converter_in_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_pixel_converter_in_endofpacket : OUT STD_LOGIC;
                    signal lcd_pixel_converter_in_ready_from_sa : OUT STD_LOGIC;
                    signal lcd_pixel_converter_in_reset_n : OUT STD_LOGIC;
                    signal lcd_pixel_converter_in_startofpacket : OUT STD_LOGIC;
                    signal lcd_pixel_converter_in_valid : OUT STD_LOGIC
                 );
end component lcd_pixel_converter_in_arbitrator;

component lcd_pixel_converter_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_in_ready_from_sa : IN STD_LOGIC;
                    signal lcd_pixel_converter_out_data : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal lcd_pixel_converter_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_pixel_converter_out_endofpacket : IN STD_LOGIC;
                    signal lcd_pixel_converter_out_startofpacket : IN STD_LOGIC;
                    signal lcd_pixel_converter_out_valid : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_pixel_converter_out_ready : OUT STD_LOGIC
                 );
end component lcd_pixel_converter_out_arbitrator;

component lcd_pixel_converter is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal empty_in : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal eop_in : IN STD_LOGIC;
                    signal ready_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sop_in : IN STD_LOGIC;
                    signal valid_in : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal empty_out : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal eop_out : OUT STD_LOGIC;
                    signal ready_out : OUT STD_LOGIC;
                    signal sop_out : OUT STD_LOGIC;
                    signal valid_out : OUT STD_LOGIC
                 );
end component lcd_pixel_converter;

component lcd_pixel_fifo_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_pixel_fifo_in_ready : IN STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_ta_sgdma_to_fifo_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_ta_sgdma_to_fifo_out_endofpacket : IN STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_out_startofpacket : IN STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_out_valid : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_pixel_fifo_in_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_pixel_fifo_in_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_pixel_fifo_in_endofpacket : OUT STD_LOGIC;
                    signal lcd_pixel_fifo_in_ready_from_sa : OUT STD_LOGIC;
                    signal lcd_pixel_fifo_in_reset_n : OUT STD_LOGIC;
                    signal lcd_pixel_fifo_in_startofpacket : OUT STD_LOGIC;
                    signal lcd_pixel_fifo_in_valid : OUT STD_LOGIC
                 );
end component lcd_pixel_fifo_in_arbitrator;

component lcd_pixel_fifo_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_pixel_fifo_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_pixel_fifo_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_pixel_fifo_out_endofpacket : IN STD_LOGIC;
                    signal lcd_pixel_fifo_out_startofpacket : IN STD_LOGIC;
                    signal lcd_pixel_fifo_out_valid : IN STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_in_ready_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_pixel_fifo_out_ready : OUT STD_LOGIC;
                    signal lcd_pixel_fifo_out_reset_n : OUT STD_LOGIC
                 );
end component lcd_pixel_fifo_out_arbitrator;

component lcd_pixel_fifo is 
           port (
                 -- inputs:
                    signal avalonst_sink_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal avalonst_sink_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal avalonst_sink_endofpacket : IN STD_LOGIC;
                    signal avalonst_sink_startofpacket : IN STD_LOGIC;
                    signal avalonst_sink_valid : IN STD_LOGIC;
                    signal avalonst_source_ready : IN STD_LOGIC;
                    signal rdclock : IN STD_LOGIC;
                    signal rdreset_n : IN STD_LOGIC;
                    signal wrclock : IN STD_LOGIC;
                    signal wrreset_n : IN STD_LOGIC;

                 -- outputs:
                    signal avalonst_sink_ready : OUT STD_LOGIC;
                    signal avalonst_source_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal avalonst_source_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal avalonst_source_endofpacket : OUT STD_LOGIC;
                    signal avalonst_source_startofpacket : OUT STD_LOGIC;
                    signal avalonst_source_valid : OUT STD_LOGIC
                 );
end component lcd_pixel_fifo;

component lcd_sgdma_csr_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_csr_irq : IN STD_LOGIC;
                    signal lcd_sgdma_csr_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr : OUT STD_LOGIC;
                    signal d1_lcd_sgdma_csr_end_xfer : OUT STD_LOGIC;
                    signal lcd_sgdma_csr_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal lcd_sgdma_csr_chipselect : OUT STD_LOGIC;
                    signal lcd_sgdma_csr_irq_from_sa : OUT STD_LOGIC;
                    signal lcd_sgdma_csr_read : OUT STD_LOGIC;
                    signal lcd_sgdma_csr_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_csr_reset_n : OUT STD_LOGIC;
                    signal lcd_sgdma_csr_write : OUT STD_LOGIC;
                    signal lcd_sgdma_csr_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component lcd_sgdma_csr_arbitrator;

component lcd_sgdma_descriptor_read_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_descriptor_read_granted_sdram_s1 : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_read : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_requests_sdram_s1 : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_sgdma_descriptor_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_descriptor_read_latency_counter : OUT STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_descriptor_read_readdatavalid : OUT STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_waitrequest : OUT STD_LOGIC
                 );
end component lcd_sgdma_descriptor_read_arbitrator;

component lcd_sgdma_descriptor_write_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_descriptor_write_granted_sdram_s1 : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_write_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_write_requests_sdram_s1 : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_write_write : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_sgdma_descriptor_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_descriptor_write_waitrequest : OUT STD_LOGIC
                 );
end component lcd_sgdma_descriptor_write_arbitrator;

component lcd_sgdma_m_read_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal lcd_sgdma_m_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_m_read_granted_sdram_s1 : IN STD_LOGIC;
                    signal lcd_sgdma_m_read_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal lcd_sgdma_m_read_read : IN STD_LOGIC;
                    signal lcd_sgdma_m_read_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal lcd_sgdma_m_read_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal lcd_sgdma_m_read_requests_sdram_s1 : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_sgdma_m_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_m_read_latency_counter : OUT STD_LOGIC;
                    signal lcd_sgdma_m_read_readdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_sgdma_m_read_readdatavalid : OUT STD_LOGIC;
                    signal lcd_sgdma_m_read_waitrequest : OUT STD_LOGIC
                 );
end component lcd_sgdma_m_read_arbitrator;

component lcd_sgdma_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_sgdma_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_sgdma_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_sgdma_out_endofpacket : IN STD_LOGIC;
                    signal lcd_sgdma_out_startofpacket : IN STD_LOGIC;
                    signal lcd_sgdma_out_valid : IN STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_in_ready_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_sgdma_out_ready : OUT STD_LOGIC
                 );
end component lcd_sgdma_out_arbitrator;

component lcd_sgdma is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal csr_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal csr_chipselect : IN STD_LOGIC;
                    signal csr_read : IN STD_LOGIC;
                    signal csr_write : IN STD_LOGIC;
                    signal csr_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_readdatavalid : IN STD_LOGIC;
                    signal descriptor_read_waitrequest : IN STD_LOGIC;
                    signal descriptor_write_waitrequest : IN STD_LOGIC;
                    signal m_read_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal m_read_readdatavalid : IN STD_LOGIC;
                    signal m_read_waitrequest : IN STD_LOGIC;
                    signal out_ready : IN STD_LOGIC;
                    signal system_reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal csr_irq : OUT STD_LOGIC;
                    signal csr_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_read : OUT STD_LOGIC;
                    signal descriptor_write_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_write_write : OUT STD_LOGIC;
                    signal descriptor_write_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m_read_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m_read_read : OUT STD_LOGIC;
                    signal out_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal out_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal out_endofpacket : OUT STD_LOGIC;
                    signal out_startofpacket : OUT STD_LOGIC;
                    signal out_valid : OUT STD_LOGIC
                 );
end component lcd_sgdma;

component lcd_sync_generator_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_out_data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal lcd_24_to_8_bits_dfa_out_empty : IN STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_out_endofpacket : IN STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_out_startofpacket : IN STD_LOGIC;
                    signal lcd_24_to_8_bits_dfa_out_valid : IN STD_LOGIC;
                    signal lcd_sync_generator_in_ready : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_sync_generator_in_data : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal lcd_sync_generator_in_empty : OUT STD_LOGIC;
                    signal lcd_sync_generator_in_endofpacket : OUT STD_LOGIC;
                    signal lcd_sync_generator_in_ready_from_sa : OUT STD_LOGIC;
                    signal lcd_sync_generator_in_reset_n : OUT STD_LOGIC;
                    signal lcd_sync_generator_in_startofpacket : OUT STD_LOGIC;
                    signal lcd_sync_generator_in_valid : OUT STD_LOGIC
                 );
end component lcd_sync_generator_in_arbitrator;

component lcd_sync_generator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal empty : IN STD_LOGIC;
                    signal eop : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sop : IN STD_LOGIC;
                    signal valid : IN STD_LOGIC;

                 -- outputs:
                    signal DEN : OUT STD_LOGIC;
                    signal HD : OUT STD_LOGIC;
                    signal RGB_OUT : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal VD : OUT STD_LOGIC;
                    signal ready : OUT STD_LOGIC
                 );
end component lcd_sync_generator;

component lcd_ta_fifo_to_dfa_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_pixel_fifo_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_pixel_fifo_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_pixel_fifo_out_endofpacket : IN STD_LOGIC;
                    signal lcd_pixel_fifo_out_startofpacket : IN STD_LOGIC;
                    signal lcd_pixel_fifo_out_valid : IN STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_in_ready : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_ta_fifo_to_dfa_in_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_ta_fifo_to_dfa_in_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_ta_fifo_to_dfa_in_endofpacket : OUT STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_in_ready_from_sa : OUT STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_in_reset_n : OUT STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_in_startofpacket : OUT STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_in_valid : OUT STD_LOGIC
                 );
end component lcd_ta_fifo_to_dfa_in_arbitrator;

component lcd_ta_fifo_to_dfa_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_64_to_32_bits_dfa_in_ready_from_sa : IN STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_ta_fifo_to_dfa_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_ta_fifo_to_dfa_out_endofpacket : IN STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_out_startofpacket : IN STD_LOGIC;
                    signal lcd_ta_fifo_to_dfa_out_valid : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_ta_fifo_to_dfa_out_ready : OUT STD_LOGIC
                 );
end component lcd_ta_fifo_to_dfa_out_arbitrator;

component lcd_ta_fifo_to_dfa is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal in_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal in_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal in_endofpacket : IN STD_LOGIC;
                    signal in_startofpacket : IN STD_LOGIC;
                    signal in_valid : IN STD_LOGIC;
                    signal out_ready : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal in_ready : OUT STD_LOGIC;
                    signal out_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal out_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal out_endofpacket : OUT STD_LOGIC;
                    signal out_startofpacket : OUT STD_LOGIC;
                    signal out_valid : OUT STD_LOGIC
                 );
end component lcd_ta_fifo_to_dfa;

component lcd_ta_sgdma_to_fifo_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_sgdma_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_sgdma_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_sgdma_out_endofpacket : IN STD_LOGIC;
                    signal lcd_sgdma_out_startofpacket : IN STD_LOGIC;
                    signal lcd_sgdma_out_valid : IN STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_in_ready : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_ta_sgdma_to_fifo_in_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_ta_sgdma_to_fifo_in_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_ta_sgdma_to_fifo_in_endofpacket : OUT STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_in_ready_from_sa : OUT STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_in_reset_n : OUT STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_in_startofpacket : OUT STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_in_valid : OUT STD_LOGIC
                 );
end component lcd_ta_sgdma_to_fifo_in_arbitrator;

component lcd_ta_sgdma_to_fifo_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_pixel_fifo_in_ready_from_sa : IN STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_out_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal lcd_ta_sgdma_to_fifo_out_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal lcd_ta_sgdma_to_fifo_out_endofpacket : IN STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_out_startofpacket : IN STD_LOGIC;
                    signal lcd_ta_sgdma_to_fifo_out_valid : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal lcd_ta_sgdma_to_fifo_out_ready : OUT STD_LOGIC
                 );
end component lcd_ta_sgdma_to_fifo_out_arbitrator;

component lcd_ta_sgdma_to_fifo is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal in_data : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal in_empty : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal in_endofpacket : IN STD_LOGIC;
                    signal in_startofpacket : IN STD_LOGIC;
                    signal in_valid : IN STD_LOGIC;
                    signal out_ready : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal in_ready : OUT STD_LOGIC;
                    signal out_data : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal out_empty : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal out_endofpacket : OUT STD_LOGIC;
                    signal out_startofpacket : OUT STD_LOGIC;
                    signal out_valid : OUT STD_LOGIC
                 );
end component lcd_ta_sgdma_to_fifo;

component performance_counter_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal performance_counter_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_granted_performance_counter_control_slave : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_performance_counter_control_slave : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_performance_counter_control_slave : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_performance_counter_control_slave : OUT STD_LOGIC;
                    signal d1_performance_counter_control_slave_end_xfer : OUT STD_LOGIC;
                    signal performance_counter_control_slave_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal performance_counter_control_slave_begintransfer : OUT STD_LOGIC;
                    signal performance_counter_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal performance_counter_control_slave_reset_n : OUT STD_LOGIC;
                    signal performance_counter_control_slave_write : OUT STD_LOGIC;
                    signal performance_counter_control_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave : OUT STD_LOGIC
                 );
end component performance_counter_control_slave_arbitrator;

component performance_counter is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal begintransfer : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component performance_counter;

component sdram_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_ddr_clock_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_descriptor_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_descriptor_read_latency_counter : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_read : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_descriptor_write_write : IN STD_LOGIC;
                    signal lcd_sgdma_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_m_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal lcd_sgdma_m_read_latency_counter : IN STD_LOGIC;
                    signal lcd_sgdma_m_read_read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal sdram_s1_readdatavalid : IN STD_LOGIC;
                    signal sdram_s1_resetrequest_n : IN STD_LOGIC;
                    signal sdram_s1_waitrequest_n : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal tse_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal tse_ddr_clock_bridge_m1_latency_counter : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal cpu_ddr_clock_bridge_m1_granted_sdram_s1 : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_ddr_clock_bridge_m1_requests_sdram_s1 : OUT STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : OUT STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_granted_sdram_s1 : OUT STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal lcd_sgdma_descriptor_read_requests_sdram_s1 : OUT STD_LOGIC;
                    signal lcd_sgdma_descriptor_write_granted_sdram_s1 : OUT STD_LOGIC;
                    signal lcd_sgdma_descriptor_write_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal lcd_sgdma_descriptor_write_requests_sdram_s1 : OUT STD_LOGIC;
                    signal lcd_sgdma_m_read_granted_sdram_s1 : OUT STD_LOGIC;
                    signal lcd_sgdma_m_read_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal lcd_sgdma_m_read_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal lcd_sgdma_m_read_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal lcd_sgdma_m_read_requests_sdram_s1 : OUT STD_LOGIC;
                    signal sdram_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal sdram_s1_beginbursttransfer : OUT STD_LOGIC;
                    signal sdram_s1_burstcount : OUT STD_LOGIC;
                    signal sdram_s1_byteenable : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal sdram_s1_read : OUT STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal sdram_s1_resetrequest_n_from_sa : OUT STD_LOGIC;
                    signal sdram_s1_waitrequest_n_from_sa : OUT STD_LOGIC;
                    signal sdram_s1_write : OUT STD_LOGIC;
                    signal sdram_s1_writedata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal tse_ddr_clock_bridge_m1_granted_sdram_s1 : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1 : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_requests_sdram_s1 : OUT STD_LOGIC
                 );
end component sdram_s1_arbitrator;

component processador_reset_clk50Mhz_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component processador_reset_clk50Mhz_domain_synch_module;

component sdram is 
           port (
                 -- inputs:
                    signal global_reset_n : IN STD_LOGIC;
                    signal local_address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal local_be : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal local_burstbegin : IN STD_LOGIC;
                    signal local_read_req : IN STD_LOGIC;
                    signal local_size : IN STD_LOGIC;
                    signal local_wdata : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal local_write_req : IN STD_LOGIC;
                    signal pll_ref_clk : IN STD_LOGIC;
                    signal soft_reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal aux_full_rate_clk : OUT STD_LOGIC;
                    signal aux_half_rate_clk : OUT STD_LOGIC;
                    signal local_init_done : OUT STD_LOGIC;
                    signal local_rdata : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal local_rdata_valid : OUT STD_LOGIC;
                    signal local_ready : OUT STD_LOGIC;
                    signal local_refresh_ack : OUT STD_LOGIC;
                    signal local_wdata_req : OUT STD_LOGIC;
                    signal mem_addr : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal mem_ba : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_cas_n : OUT STD_LOGIC;
                    signal mem_cke : OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
                    signal mem_clk : INOUT STD_LOGIC_VECTOR (0 DOWNTO 0);
                    signal mem_clk_n : INOUT STD_LOGIC_VECTOR (0 DOWNTO 0);
                    signal mem_cs_n : OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
                    signal mem_dm : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_dq : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal mem_dqs : INOUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_ras_n : OUT STD_LOGIC;
                    signal mem_we_n : OUT STD_LOGIC;
                    signal phy_clk : OUT STD_LOGIC;
                    signal reset_phy_clk_n : OUT STD_LOGIC;
                    signal reset_request_n : OUT STD_LOGIC
                 );
end component sdram;

component sgdma_rx_csr_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_csr_irq : IN STD_LOGIC;
                    signal sgdma_rx_csr_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal cpuNios_data_master_granted_sgdma_rx_csr : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_sgdma_rx_csr : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_sgdma_rx_csr : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_sgdma_rx_csr : OUT STD_LOGIC;
                    signal d1_sgdma_rx_csr_end_xfer : OUT STD_LOGIC;
                    signal sgdma_rx_csr_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal sgdma_rx_csr_chipselect : OUT STD_LOGIC;
                    signal sgdma_rx_csr_irq_from_sa : OUT STD_LOGIC;
                    signal sgdma_rx_csr_read : OUT STD_LOGIC;
                    signal sgdma_rx_csr_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_csr_reset_n : OUT STD_LOGIC;
                    signal sgdma_rx_csr_write : OUT STD_LOGIC;
                    signal sgdma_rx_csr_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sgdma_rx_csr_arbitrator;

component sgdma_rx_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_in_ready : IN STD_LOGIC;
                    signal tse_mac_receive_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_receive_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal tse_mac_receive_endofpacket : IN STD_LOGIC;
                    signal tse_mac_receive_error : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal tse_mac_receive_startofpacket : IN STD_LOGIC;
                    signal tse_mac_receive_valid : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_rx_in_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_in_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sgdma_rx_in_endofpacket : OUT STD_LOGIC;
                    signal sgdma_rx_in_error : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal sgdma_rx_in_ready_from_sa : OUT STD_LOGIC;
                    signal sgdma_rx_in_startofpacket : OUT STD_LOGIC;
                    signal sgdma_rx_in_valid : OUT STD_LOGIC
                 );
end component sgdma_rx_in_arbitrator;

component sgdma_rx_descriptor_read_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_descriptor_offset_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal descriptor_offset_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (255 DOWNTO 0);
                    signal descriptor_offset_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_read : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_rx_descriptor_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_read_latency_counter : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_read_readdatavalid : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_rx_descriptor_read_arbitrator;

component sgdma_rx_descriptor_write_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_descriptor_offset_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal descriptor_offset_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_write : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal sgdma_rx_descriptor_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_write_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_rx_descriptor_write_arbitrator;

component sgdma_rx_m_write_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_tse_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_m_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_write : IN STD_LOGIC;
                    signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_rx_m_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_m_write_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_rx_m_write_arbitrator;

component sgdma_rx is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal csr_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal csr_chipselect : IN STD_LOGIC;
                    signal csr_read : IN STD_LOGIC;
                    signal csr_write : IN STD_LOGIC;
                    signal csr_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_readdatavalid : IN STD_LOGIC;
                    signal descriptor_read_waitrequest : IN STD_LOGIC;
                    signal descriptor_write_waitrequest : IN STD_LOGIC;
                    signal in_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal in_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal in_endofpacket : IN STD_LOGIC;
                    signal in_error : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal in_startofpacket : IN STD_LOGIC;
                    signal in_valid : IN STD_LOGIC;
                    signal m_write_waitrequest : IN STD_LOGIC;
                    signal system_reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal csr_irq : OUT STD_LOGIC;
                    signal csr_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_read : OUT STD_LOGIC;
                    signal descriptor_write_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_write_write : OUT STD_LOGIC;
                    signal descriptor_write_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal in_ready : OUT STD_LOGIC;
                    signal m_write_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m_write_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_write_write : OUT STD_LOGIC;
                    signal m_write_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sgdma_rx;

component sgdma_tx_csr_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_csr_irq : IN STD_LOGIC;
                    signal sgdma_tx_csr_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal cpuNios_data_master_granted_sgdma_tx_csr : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_sgdma_tx_csr : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_sgdma_tx_csr : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_sgdma_tx_csr : OUT STD_LOGIC;
                    signal d1_sgdma_tx_csr_end_xfer : OUT STD_LOGIC;
                    signal sgdma_tx_csr_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal sgdma_tx_csr_chipselect : OUT STD_LOGIC;
                    signal sgdma_tx_csr_irq_from_sa : OUT STD_LOGIC;
                    signal sgdma_tx_csr_read : OUT STD_LOGIC;
                    signal sgdma_tx_csr_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_csr_reset_n : OUT STD_LOGIC;
                    signal sgdma_tx_csr_write : OUT STD_LOGIC;
                    signal sgdma_tx_csr_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sgdma_tx_csr_arbitrator;

component sgdma_tx_descriptor_read_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_descriptor_offset_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal descriptor_offset_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (255 DOWNTO 0);
                    signal descriptor_offset_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_read : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_tx_descriptor_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_read_latency_counter : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_read_readdatavalid : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_tx_descriptor_read_arbitrator;

component sgdma_tx_descriptor_write_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_descriptor_offset_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal descriptor_offset_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_write : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal sgdma_tx_descriptor_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_write_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_tx_descriptor_write_arbitrator;

component sgdma_tx_m_read_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_tse_ddr_clock_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_m_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1_shift_register : IN STD_LOGIC;
                    signal sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_ddr_clock_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_tx_m_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_latency_counter : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_readdatavalid : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_tx_m_read_arbitrator;

component sgdma_tx_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sgdma_tx_out_endofpacket : IN STD_LOGIC;
                    signal sgdma_tx_out_error : IN STD_LOGIC;
                    signal sgdma_tx_out_startofpacket : IN STD_LOGIC;
                    signal sgdma_tx_out_valid : IN STD_LOGIC;
                    signal tse_mac_transmit_ready_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_tx_out_ready : OUT STD_LOGIC
                 );
end component sgdma_tx_out_arbitrator;

component sgdma_tx is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal csr_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal csr_chipselect : IN STD_LOGIC;
                    signal csr_read : IN STD_LOGIC;
                    signal csr_write : IN STD_LOGIC;
                    signal csr_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_readdatavalid : IN STD_LOGIC;
                    signal descriptor_read_waitrequest : IN STD_LOGIC;
                    signal descriptor_write_waitrequest : IN STD_LOGIC;
                    signal m_read_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m_read_readdatavalid : IN STD_LOGIC;
                    signal m_read_waitrequest : IN STD_LOGIC;
                    signal out_ready : IN STD_LOGIC;
                    signal system_reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal csr_irq : OUT STD_LOGIC;
                    signal csr_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_read : OUT STD_LOGIC;
                    signal descriptor_write_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_write_write : OUT STD_LOGIC;
                    signal descriptor_write_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m_read_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m_read_read : OUT STD_LOGIC;
                    signal out_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal out_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal out_endofpacket : OUT STD_LOGIC;
                    signal out_error : OUT STD_LOGIC;
                    signal out_startofpacket : OUT STD_LOGIC;
                    signal out_valid : OUT STD_LOGIC
                 );
end component sgdma_tx;

component sys_clk_timer_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_timer_s1_irq : IN STD_LOGIC;
                    signal sys_clk_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal cpuNios_data_master_granted_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal d1_sys_clk_timer_s1_end_xfer : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal sys_clk_timer_s1_chipselect : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_irq_from_sa : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sys_clk_timer_s1_reset_n : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_write_n : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sys_clk_timer_s1_arbitrator;

component sys_clk_timer is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sys_clk_timer;

component sysid_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal cpuNios_data_master_granted_sysid_control_slave : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_sysid_control_slave : OUT STD_LOGIC;
                    signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                    signal sysid_control_slave_address : OUT STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sysid_control_slave_reset_n : OUT STD_LOGIC
                 );
end component sysid_control_slave_arbitrator;

component sysid is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC;
                    signal clock : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sysid;

component tse_ddr_clock_bridge_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_m_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal sgdma_rx_m_write_write : IN STD_LOGIC;
                    signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_latency_counter : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_s1_endofpacket : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_ddr_clock_bridge_s1_readdatavalid : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_s1_waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal d1_tse_ddr_clock_bridge_s1_end_xfer : OUT STD_LOGIC;
                    signal sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal tse_ddr_clock_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal tse_ddr_clock_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal tse_ddr_clock_bridge_s1_read : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_ddr_clock_bridge_s1_reset_n : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_s1_write : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component tse_ddr_clock_bridge_s1_arbitrator;

component tse_ddr_clock_bridge_m1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_sdram_s1_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
                    signal sdram_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal tse_ddr_clock_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal tse_ddr_clock_bridge_m1_granted_sdram_s1 : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_read : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1 : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_requests_sdram_s1 : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_write : IN STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal tse_ddr_clock_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal tse_ddr_clock_bridge_m1_latency_counter : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_ddr_clock_bridge_m1_readdatavalid : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_reset_n : OUT STD_LOGIC;
                    signal tse_ddr_clock_bridge_m1_waitrequest : OUT STD_LOGIC
                 );
end component tse_ddr_clock_bridge_m1_arbitrator;

component tse_ddr_clock_bridge is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_readdatavalid : IN STD_LOGIC;
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_readdatavalid : OUT STD_LOGIC;
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component tse_ddr_clock_bridge;

component tse_ddr_clock_bridge_bridge_arbitrator is 
end component tse_ddr_clock_bridge_bridge_arbitrator;

component tse_mac_control_port_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpuNios_data_master_address_to_slave : IN STD_LOGIC_VECTOR (26 DOWNTO 0);
                    signal cpuNios_data_master_read : IN STD_LOGIC;
                    signal cpuNios_data_master_waitrequest : IN STD_LOGIC;
                    signal cpuNios_data_master_write : IN STD_LOGIC;
                    signal cpuNios_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal tse_mac_control_port_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_control_port_waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal cpuNios_data_master_granted_tse_mac_control_port : OUT STD_LOGIC;
                    signal cpuNios_data_master_qualified_request_tse_mac_control_port : OUT STD_LOGIC;
                    signal cpuNios_data_master_read_data_valid_tse_mac_control_port : OUT STD_LOGIC;
                    signal cpuNios_data_master_requests_tse_mac_control_port : OUT STD_LOGIC;
                    signal d1_tse_mac_control_port_end_xfer : OUT STD_LOGIC;
                    signal tse_mac_control_port_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal tse_mac_control_port_read : OUT STD_LOGIC;
                    signal tse_mac_control_port_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_control_port_reset : OUT STD_LOGIC;
                    signal tse_mac_control_port_waitrequest_from_sa : OUT STD_LOGIC;
                    signal tse_mac_control_port_write : OUT STD_LOGIC;
                    signal tse_mac_control_port_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component tse_mac_control_port_arbitrator;

component tse_mac_transmit_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sgdma_tx_out_endofpacket : IN STD_LOGIC;
                    signal sgdma_tx_out_error : IN STD_LOGIC;
                    signal sgdma_tx_out_startofpacket : IN STD_LOGIC;
                    signal sgdma_tx_out_valid : IN STD_LOGIC;
                    signal tse_mac_transmit_ready : IN STD_LOGIC;

                 -- outputs:
                    signal tse_mac_transmit_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_transmit_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal tse_mac_transmit_endofpacket : OUT STD_LOGIC;
                    signal tse_mac_transmit_error : OUT STD_LOGIC;
                    signal tse_mac_transmit_ready_from_sa : OUT STD_LOGIC;
                    signal tse_mac_transmit_startofpacket : OUT STD_LOGIC;
                    signal tse_mac_transmit_valid : OUT STD_LOGIC
                 );
end component tse_mac_transmit_arbitrator;

component tse_mac_receive_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_in_ready_from_sa : IN STD_LOGIC;
                    signal tse_mac_receive_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_receive_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal tse_mac_receive_endofpacket : IN STD_LOGIC;
                    signal tse_mac_receive_error : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal tse_mac_receive_startofpacket : IN STD_LOGIC;
                    signal tse_mac_receive_valid : IN STD_LOGIC;

                 -- outputs:
                    signal tse_mac_receive_ready : OUT STD_LOGIC
                 );
end component tse_mac_receive_arbitrator;

component tse_mac is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal ff_rx_clk : IN STD_LOGIC;
                    signal ff_rx_rdy : IN STD_LOGIC;
                    signal ff_tx_clk : IN STD_LOGIC;
                    signal ff_tx_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ff_tx_eop : IN STD_LOGIC;
                    signal ff_tx_err : IN STD_LOGIC;
                    signal ff_tx_mod : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ff_tx_sop : IN STD_LOGIC;
                    signal ff_tx_wren : IN STD_LOGIC;
                    signal gm_rx_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_rx_dv : IN STD_LOGIC;
                    signal gm_rx_err : IN STD_LOGIC;
                    signal m_rx_col : IN STD_LOGIC;
                    signal m_rx_crs : IN STD_LOGIC;
                    signal m_rx_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_rx_en : IN STD_LOGIC;
                    signal m_rx_err : IN STD_LOGIC;
                    signal mdio_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal rx_clk : IN STD_LOGIC;
                    signal set_10 : IN STD_LOGIC;
                    signal set_1000 : IN STD_LOGIC;
                    signal tx_clk : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal ena_10 : OUT STD_LOGIC;
                    signal eth_mode : OUT STD_LOGIC;
                    signal ff_rx_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ff_rx_dval : OUT STD_LOGIC;
                    signal ff_rx_eop : OUT STD_LOGIC;
                    signal ff_rx_mod : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ff_rx_sop : OUT STD_LOGIC;
                    signal ff_tx_rdy : OUT STD_LOGIC;
                    signal gm_tx_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_tx_en : OUT STD_LOGIC;
                    signal gm_tx_err : OUT STD_LOGIC;
                    signal m_tx_d : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_tx_en : OUT STD_LOGIC;
                    signal m_tx_err : OUT STD_LOGIC;
                    signal mdc : OUT STD_LOGIC;
                    signal mdio_oen : OUT STD_LOGIC;
                    signal mdio_out : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal rx_err : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal waitrequest : OUT STD_LOGIC
                 );
end component tse_mac;

component processador_reset_clk100MHz_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component processador_reset_clk100MHz_domain_synch_module;

component processador_reset_sdram_phy_clk_out_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component processador_reset_sdram_phy_clk_out_domain_synch_module;

                signal clk100MHz_reset_n :  STD_LOGIC;
                signal clk50Mhz_reset_n :  STD_LOGIC;
                signal cpuNios_data_master_address :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal cpuNios_data_master_address_to_slave :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal cpuNios_data_master_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpuNios_data_master_debugaccess :  STD_LOGIC;
                signal cpuNios_data_master_granted_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_data_master_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 :  STD_LOGIC;
                signal cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal cpuNios_data_master_granted_lcd_i2c_en_s1 :  STD_LOGIC;
                signal cpuNios_data_master_granted_lcd_i2c_scl_s1 :  STD_LOGIC;
                signal cpuNios_data_master_granted_lcd_i2c_sdat_s1 :  STD_LOGIC;
                signal cpuNios_data_master_granted_performance_counter_control_slave :  STD_LOGIC;
                signal cpuNios_data_master_granted_sgdma_rx_csr :  STD_LOGIC;
                signal cpuNios_data_master_granted_sgdma_tx_csr :  STD_LOGIC;
                signal cpuNios_data_master_granted_sys_clk_timer_s1 :  STD_LOGIC;
                signal cpuNios_data_master_granted_sysid_control_slave :  STD_LOGIC;
                signal cpuNios_data_master_granted_tse_mac_control_port :  STD_LOGIC;
                signal cpuNios_data_master_irq :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_lcd_i2c_en_s1 :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_performance_counter_control_slave :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_sgdma_rx_csr :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_sgdma_tx_csr :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_sys_clk_timer_s1 :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal cpuNios_data_master_qualified_request_tse_mac_control_port :  STD_LOGIC;
                signal cpuNios_data_master_read :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_descriptor_memory_s1 :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_fft_pipeline_0_avalon_slave_0 :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_lcd_i2c_en_s1 :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_lcd_i2c_scl_s1 :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_lcd_i2c_sdat_s1 :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_performance_counter_control_slave :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_sgdma_rx_csr :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_sgdma_tx_csr :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_sys_clk_timer_s1 :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_sysid_control_slave :  STD_LOGIC;
                signal cpuNios_data_master_read_data_valid_tse_mac_control_port :  STD_LOGIC;
                signal cpuNios_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpuNios_data_master_requests_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_data_master_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 :  STD_LOGIC;
                signal cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal cpuNios_data_master_requests_lcd_i2c_en_s1 :  STD_LOGIC;
                signal cpuNios_data_master_requests_lcd_i2c_scl_s1 :  STD_LOGIC;
                signal cpuNios_data_master_requests_lcd_i2c_sdat_s1 :  STD_LOGIC;
                signal cpuNios_data_master_requests_performance_counter_control_slave :  STD_LOGIC;
                signal cpuNios_data_master_requests_sgdma_rx_csr :  STD_LOGIC;
                signal cpuNios_data_master_requests_sgdma_tx_csr :  STD_LOGIC;
                signal cpuNios_data_master_requests_sys_clk_timer_s1 :  STD_LOGIC;
                signal cpuNios_data_master_requests_sysid_control_slave :  STD_LOGIC;
                signal cpuNios_data_master_requests_tse_mac_control_port :  STD_LOGIC;
                signal cpuNios_data_master_waitrequest :  STD_LOGIC;
                signal cpuNios_data_master_write :  STD_LOGIC;
                signal cpuNios_data_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpuNios_instruction_master_address :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal cpuNios_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal cpuNios_instruction_master_granted_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_instruction_master_read :  STD_LOGIC;
                signal cpuNios_instruction_master_read_data_valid_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register :  STD_LOGIC;
                signal cpuNios_instruction_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpuNios_instruction_master_requests_cpuNios_jtag_debug_module :  STD_LOGIC;
                signal cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal cpuNios_instruction_master_waitrequest :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal cpuNios_jtag_debug_module_begintransfer :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpuNios_jtag_debug_module_chipselect :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_debugaccess :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpuNios_jtag_debug_module_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpuNios_jtag_debug_module_reset_n :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_resetrequest :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_resetrequest_from_sa :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_write :  STD_LOGIC;
                signal cpuNios_jtag_debug_module_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_address :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_endofpacket :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_granted_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_latency_counter :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_nativeaddress :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_read :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_readdatavalid :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_requests_sdram_s1 :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_reset_n :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_waitrequest :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_write :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_endofpacket :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_nativeaddress :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_read :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_readdatavalid :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_reset_n :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_waitrequest :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_write :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal d1_cpuNios_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal d1_cpu_ddr_clock_bridge_s1_end_xfer :  STD_LOGIC;
                signal d1_descriptor_memory_s1_end_xfer :  STD_LOGIC;
                signal d1_descriptor_offset_bridge_s1_end_xfer :  STD_LOGIC;
                signal d1_fft_pipeline_0_avalon_slave_0_end_xfer :  STD_LOGIC;
                signal d1_jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal d1_lcd_i2c_en_s1_end_xfer :  STD_LOGIC;
                signal d1_lcd_i2c_scl_s1_end_xfer :  STD_LOGIC;
                signal d1_lcd_i2c_sdat_s1_end_xfer :  STD_LOGIC;
                signal d1_lcd_sgdma_csr_end_xfer :  STD_LOGIC;
                signal d1_performance_counter_control_slave_end_xfer :  STD_LOGIC;
                signal d1_sdram_s1_end_xfer :  STD_LOGIC;
                signal d1_sgdma_rx_csr_end_xfer :  STD_LOGIC;
                signal d1_sgdma_tx_csr_end_xfer :  STD_LOGIC;
                signal d1_sys_clk_timer_s1_end_xfer :  STD_LOGIC;
                signal d1_sysid_control_slave_end_xfer :  STD_LOGIC;
                signal d1_tse_ddr_clock_bridge_s1_end_xfer :  STD_LOGIC;
                signal d1_tse_mac_control_port_end_xfer :  STD_LOGIC;
                signal descriptor_memory_s1_address :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal descriptor_memory_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_memory_s1_chipselect :  STD_LOGIC;
                signal descriptor_memory_s1_clken :  STD_LOGIC;
                signal descriptor_memory_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal descriptor_memory_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal descriptor_memory_s1_reset :  STD_LOGIC;
                signal descriptor_memory_s1_write :  STD_LOGIC;
                signal descriptor_memory_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal descriptor_offset_bridge_m1_address :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal descriptor_offset_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (26 DOWNTO 0);
                signal descriptor_offset_bridge_m1_burstcount :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_byteenable :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_offset_bridge_m1_chipselect :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_dbs_address :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_offset_bridge_m1_dbs_write_32 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal descriptor_offset_bridge_m1_debugaccess :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_endofpacket :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_latency_counter :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_read :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1 :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_readdata :  STD_LOGIC_VECTOR (255 DOWNTO 0);
                signal descriptor_offset_bridge_m1_readdatavalid :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_waitrequest :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_write :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_writedata :  STD_LOGIC_VECTOR (255 DOWNTO 0);
                signal descriptor_offset_bridge_s1_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal descriptor_offset_bridge_s1_arbiterlock :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_arbiterlock2 :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_burstcount :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_byteenable :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal descriptor_offset_bridge_s1_chipselect :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_debugaccess :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_endofpacket :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_nativeaddress :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal descriptor_offset_bridge_s1_read :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_readdata :  STD_LOGIC_VECTOR (255 DOWNTO 0);
                signal descriptor_offset_bridge_s1_readdata_from_sa :  STD_LOGIC_VECTOR (255 DOWNTO 0);
                signal descriptor_offset_bridge_s1_readdatavalid :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_reset_n :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_waitrequest :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_write :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_writedata :  STD_LOGIC_VECTOR (255 DOWNTO 0);
                signal fft_pipeline_0_avalon_slave_0_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal fft_pipeline_0_avalon_slave_0_chipselect :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal fft_pipeline_0_avalon_slave_0_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal fft_pipeline_0_avalon_slave_0_reset :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_write :  STD_LOGIC;
                signal fft_pipeline_0_avalon_slave_0_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_DEN_from_the_lcd_sync_generator :  STD_LOGIC;
                signal internal_HD_from_the_lcd_sync_generator :  STD_LOGIC;
                signal internal_RGB_OUT_from_the_lcd_sync_generator :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_VD_from_the_lcd_sync_generator :  STD_LOGIC;
                signal internal_counter_from_the_fft_pipeline_0 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal internal_ena_10_from_the_tse_mac :  STD_LOGIC;
                signal internal_eth_mode_from_the_tse_mac :  STD_LOGIC;
                signal internal_gm_tx_d_from_the_tse_mac :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_gm_tx_en_from_the_tse_mac :  STD_LOGIC;
                signal internal_gm_tx_err_from_the_tse_mac :  STD_LOGIC;
                signal internal_local_init_done_from_the_sdram :  STD_LOGIC;
                signal internal_local_refresh_ack_from_the_sdram :  STD_LOGIC;
                signal internal_local_wdata_req_from_the_sdram :  STD_LOGIC;
                signal internal_m_tx_d_from_the_tse_mac :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_m_tx_en_from_the_tse_mac :  STD_LOGIC;
                signal internal_m_tx_err_from_the_tse_mac :  STD_LOGIC;
                signal internal_mdc_from_the_tse_mac :  STD_LOGIC;
                signal internal_mdio_oen_from_the_tse_mac :  STD_LOGIC;
                signal internal_mdio_out_from_the_tse_mac :  STD_LOGIC;
                signal internal_mem_addr_from_the_sdram :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal internal_mem_ba_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_mem_cas_n_from_the_sdram :  STD_LOGIC;
                signal internal_mem_cke_from_the_sdram :  STD_LOGIC;
                signal internal_mem_cs_n_from_the_sdram :  STD_LOGIC;
                signal internal_mem_dm_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_mem_ras_n_from_the_sdram :  STD_LOGIC;
                signal internal_mem_we_n_from_the_sdram :  STD_LOGIC;
                signal internal_out_port_from_the_lcd_i2c_en :  STD_LOGIC;
                signal internal_out_port_from_the_lcd_i2c_scl :  STD_LOGIC;
                signal internal_reset_phy_clk_n_from_the_sdram :  STD_LOGIC;
                signal internal_sdram_phy_clk_out :  STD_LOGIC;
                signal internal_tx_out_from_the_fft_pipeline_0 :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_address :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_chipselect :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_read_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readyfordata :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reset_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_write_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_24_to_8_bits_dfa_in_data :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal lcd_24_to_8_bits_dfa_in_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal lcd_24_to_8_bits_dfa_in_endofpacket :  STD_LOGIC;
                signal lcd_24_to_8_bits_dfa_in_ready :  STD_LOGIC;
                signal lcd_24_to_8_bits_dfa_in_ready_from_sa :  STD_LOGIC;
                signal lcd_24_to_8_bits_dfa_in_reset_n :  STD_LOGIC;
                signal lcd_24_to_8_bits_dfa_in_startofpacket :  STD_LOGIC;
                signal lcd_24_to_8_bits_dfa_in_valid :  STD_LOGIC;
                signal lcd_24_to_8_bits_dfa_out_data :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal lcd_24_to_8_bits_dfa_out_empty :  STD_LOGIC;
                signal lcd_24_to_8_bits_dfa_out_endofpacket :  STD_LOGIC;
                signal lcd_24_to_8_bits_dfa_out_ready :  STD_LOGIC;
                signal lcd_24_to_8_bits_dfa_out_startofpacket :  STD_LOGIC;
                signal lcd_24_to_8_bits_dfa_out_valid :  STD_LOGIC;
                signal lcd_64_to_32_bits_dfa_in_data :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal lcd_64_to_32_bits_dfa_in_empty :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_64_to_32_bits_dfa_in_endofpacket :  STD_LOGIC;
                signal lcd_64_to_32_bits_dfa_in_ready :  STD_LOGIC;
                signal lcd_64_to_32_bits_dfa_in_ready_from_sa :  STD_LOGIC;
                signal lcd_64_to_32_bits_dfa_in_reset_n :  STD_LOGIC;
                signal lcd_64_to_32_bits_dfa_in_startofpacket :  STD_LOGIC;
                signal lcd_64_to_32_bits_dfa_in_valid :  STD_LOGIC;
                signal lcd_64_to_32_bits_dfa_out_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_64_to_32_bits_dfa_out_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal lcd_64_to_32_bits_dfa_out_endofpacket :  STD_LOGIC;
                signal lcd_64_to_32_bits_dfa_out_ready :  STD_LOGIC;
                signal lcd_64_to_32_bits_dfa_out_startofpacket :  STD_LOGIC;
                signal lcd_64_to_32_bits_dfa_out_valid :  STD_LOGIC;
                signal lcd_i2c_en_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal lcd_i2c_en_s1_chipselect :  STD_LOGIC;
                signal lcd_i2c_en_s1_readdata :  STD_LOGIC;
                signal lcd_i2c_en_s1_readdata_from_sa :  STD_LOGIC;
                signal lcd_i2c_en_s1_reset_n :  STD_LOGIC;
                signal lcd_i2c_en_s1_write_n :  STD_LOGIC;
                signal lcd_i2c_en_s1_writedata :  STD_LOGIC;
                signal lcd_i2c_scl_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal lcd_i2c_scl_s1_chipselect :  STD_LOGIC;
                signal lcd_i2c_scl_s1_readdata :  STD_LOGIC;
                signal lcd_i2c_scl_s1_readdata_from_sa :  STD_LOGIC;
                signal lcd_i2c_scl_s1_reset_n :  STD_LOGIC;
                signal lcd_i2c_scl_s1_write_n :  STD_LOGIC;
                signal lcd_i2c_scl_s1_writedata :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal lcd_i2c_sdat_s1_chipselect :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_readdata :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_readdata_from_sa :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_reset_n :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_write_n :  STD_LOGIC;
                signal lcd_i2c_sdat_s1_writedata :  STD_LOGIC;
                signal lcd_pixel_converter_in_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_pixel_converter_in_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal lcd_pixel_converter_in_endofpacket :  STD_LOGIC;
                signal lcd_pixel_converter_in_ready :  STD_LOGIC;
                signal lcd_pixel_converter_in_ready_from_sa :  STD_LOGIC;
                signal lcd_pixel_converter_in_reset_n :  STD_LOGIC;
                signal lcd_pixel_converter_in_startofpacket :  STD_LOGIC;
                signal lcd_pixel_converter_in_valid :  STD_LOGIC;
                signal lcd_pixel_converter_out_data :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal lcd_pixel_converter_out_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal lcd_pixel_converter_out_endofpacket :  STD_LOGIC;
                signal lcd_pixel_converter_out_ready :  STD_LOGIC;
                signal lcd_pixel_converter_out_startofpacket :  STD_LOGIC;
                signal lcd_pixel_converter_out_valid :  STD_LOGIC;
                signal lcd_pixel_fifo_in_data :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal lcd_pixel_fifo_in_empty :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_pixel_fifo_in_endofpacket :  STD_LOGIC;
                signal lcd_pixel_fifo_in_ready :  STD_LOGIC;
                signal lcd_pixel_fifo_in_ready_from_sa :  STD_LOGIC;
                signal lcd_pixel_fifo_in_reset_n :  STD_LOGIC;
                signal lcd_pixel_fifo_in_startofpacket :  STD_LOGIC;
                signal lcd_pixel_fifo_in_valid :  STD_LOGIC;
                signal lcd_pixel_fifo_out_data :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal lcd_pixel_fifo_out_empty :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_pixel_fifo_out_endofpacket :  STD_LOGIC;
                signal lcd_pixel_fifo_out_ready :  STD_LOGIC;
                signal lcd_pixel_fifo_out_reset_n :  STD_LOGIC;
                signal lcd_pixel_fifo_out_startofpacket :  STD_LOGIC;
                signal lcd_pixel_fifo_out_valid :  STD_LOGIC;
                signal lcd_sgdma_csr_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal lcd_sgdma_csr_chipselect :  STD_LOGIC;
                signal lcd_sgdma_csr_irq :  STD_LOGIC;
                signal lcd_sgdma_csr_irq_from_sa :  STD_LOGIC;
                signal lcd_sgdma_csr_read :  STD_LOGIC;
                signal lcd_sgdma_csr_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_csr_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_csr_reset_n :  STD_LOGIC;
                signal lcd_sgdma_csr_write :  STD_LOGIC;
                signal lcd_sgdma_csr_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_descriptor_read_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_descriptor_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_descriptor_read_granted_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_latency_counter :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_qualified_request_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_read :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_descriptor_read_readdatavalid :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_requests_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_read_waitrequest :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_descriptor_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_descriptor_write_granted_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_qualified_request_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_requests_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_waitrequest :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_write :  STD_LOGIC;
                signal lcd_sgdma_descriptor_write_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_m_read_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_m_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_sgdma_m_read_granted_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_m_read_latency_counter :  STD_LOGIC;
                signal lcd_sgdma_m_read_qualified_request_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_m_read_read :  STD_LOGIC;
                signal lcd_sgdma_m_read_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_m_read_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal lcd_sgdma_m_read_readdata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal lcd_sgdma_m_read_readdatavalid :  STD_LOGIC;
                signal lcd_sgdma_m_read_requests_sdram_s1 :  STD_LOGIC;
                signal lcd_sgdma_m_read_waitrequest :  STD_LOGIC;
                signal lcd_sgdma_out_data :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal lcd_sgdma_out_empty :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_sgdma_out_endofpacket :  STD_LOGIC;
                signal lcd_sgdma_out_ready :  STD_LOGIC;
                signal lcd_sgdma_out_startofpacket :  STD_LOGIC;
                signal lcd_sgdma_out_valid :  STD_LOGIC;
                signal lcd_sync_generator_in_data :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal lcd_sync_generator_in_empty :  STD_LOGIC;
                signal lcd_sync_generator_in_endofpacket :  STD_LOGIC;
                signal lcd_sync_generator_in_ready :  STD_LOGIC;
                signal lcd_sync_generator_in_ready_from_sa :  STD_LOGIC;
                signal lcd_sync_generator_in_reset_n :  STD_LOGIC;
                signal lcd_sync_generator_in_startofpacket :  STD_LOGIC;
                signal lcd_sync_generator_in_valid :  STD_LOGIC;
                signal lcd_ta_fifo_to_dfa_in_data :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal lcd_ta_fifo_to_dfa_in_empty :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_ta_fifo_to_dfa_in_endofpacket :  STD_LOGIC;
                signal lcd_ta_fifo_to_dfa_in_ready :  STD_LOGIC;
                signal lcd_ta_fifo_to_dfa_in_ready_from_sa :  STD_LOGIC;
                signal lcd_ta_fifo_to_dfa_in_reset_n :  STD_LOGIC;
                signal lcd_ta_fifo_to_dfa_in_startofpacket :  STD_LOGIC;
                signal lcd_ta_fifo_to_dfa_in_valid :  STD_LOGIC;
                signal lcd_ta_fifo_to_dfa_out_data :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal lcd_ta_fifo_to_dfa_out_empty :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_ta_fifo_to_dfa_out_endofpacket :  STD_LOGIC;
                signal lcd_ta_fifo_to_dfa_out_ready :  STD_LOGIC;
                signal lcd_ta_fifo_to_dfa_out_startofpacket :  STD_LOGIC;
                signal lcd_ta_fifo_to_dfa_out_valid :  STD_LOGIC;
                signal lcd_ta_sgdma_to_fifo_in_data :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal lcd_ta_sgdma_to_fifo_in_empty :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_ta_sgdma_to_fifo_in_endofpacket :  STD_LOGIC;
                signal lcd_ta_sgdma_to_fifo_in_ready :  STD_LOGIC;
                signal lcd_ta_sgdma_to_fifo_in_ready_from_sa :  STD_LOGIC;
                signal lcd_ta_sgdma_to_fifo_in_reset_n :  STD_LOGIC;
                signal lcd_ta_sgdma_to_fifo_in_startofpacket :  STD_LOGIC;
                signal lcd_ta_sgdma_to_fifo_in_valid :  STD_LOGIC;
                signal lcd_ta_sgdma_to_fifo_out_data :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal lcd_ta_sgdma_to_fifo_out_empty :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_ta_sgdma_to_fifo_out_endofpacket :  STD_LOGIC;
                signal lcd_ta_sgdma_to_fifo_out_ready :  STD_LOGIC;
                signal lcd_ta_sgdma_to_fifo_out_startofpacket :  STD_LOGIC;
                signal lcd_ta_sgdma_to_fifo_out_valid :  STD_LOGIC;
                signal module_input30 :  STD_LOGIC;
                signal module_input43 :  STD_LOGIC;
                signal module_input44 :  STD_LOGIC;
                signal out_clk_sdram_aux_full_rate_clk :  STD_LOGIC;
                signal out_clk_sdram_aux_half_rate_clk :  STD_LOGIC;
                signal out_clk_sdram_phy_clk :  STD_LOGIC;
                signal performance_counter_control_slave_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal performance_counter_control_slave_begintransfer :  STD_LOGIC;
                signal performance_counter_control_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal performance_counter_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal performance_counter_control_slave_reset_n :  STD_LOGIC;
                signal performance_counter_control_slave_write :  STD_LOGIC;
                signal performance_counter_control_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1 :  STD_LOGIC;
                signal registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave :  STD_LOGIC;
                signal reset_n_sources :  STD_LOGIC;
                signal sdram_phy_clk_out_reset_n :  STD_LOGIC;
                signal sdram_s1_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal sdram_s1_beginbursttransfer :  STD_LOGIC;
                signal sdram_s1_burstcount :  STD_LOGIC;
                signal sdram_s1_byteenable :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal sdram_s1_read :  STD_LOGIC;
                signal sdram_s1_readdata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal sdram_s1_readdata_from_sa :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal sdram_s1_readdatavalid :  STD_LOGIC;
                signal sdram_s1_resetrequest_n :  STD_LOGIC;
                signal sdram_s1_resetrequest_n_from_sa :  STD_LOGIC;
                signal sdram_s1_waitrequest_n :  STD_LOGIC;
                signal sdram_s1_waitrequest_n_from_sa :  STD_LOGIC;
                signal sdram_s1_write :  STD_LOGIC;
                signal sdram_s1_writedata :  STD_LOGIC_VECTOR (63 DOWNTO 0);
                signal sgdma_rx_csr_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sgdma_rx_csr_chipselect :  STD_LOGIC;
                signal sgdma_rx_csr_irq :  STD_LOGIC;
                signal sgdma_rx_csr_irq_from_sa :  STD_LOGIC;
                signal sgdma_rx_csr_read :  STD_LOGIC;
                signal sgdma_rx_csr_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_csr_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_csr_reset_n :  STD_LOGIC;
                signal sgdma_rx_csr_write :  STD_LOGIC;
                signal sgdma_rx_csr_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_read_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_latency_counter :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_read_readdatavalid :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_waitrequest :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_waitrequest :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_write :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_in_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_in_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sgdma_rx_in_endofpacket :  STD_LOGIC;
                signal sgdma_rx_in_error :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal sgdma_rx_in_ready :  STD_LOGIC;
                signal sgdma_rx_in_ready_from_sa :  STD_LOGIC;
                signal sgdma_rx_in_startofpacket :  STD_LOGIC;
                signal sgdma_rx_in_valid :  STD_LOGIC;
                signal sgdma_rx_m_write_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_m_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_m_write_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal sgdma_rx_m_write_waitrequest :  STD_LOGIC;
                signal sgdma_rx_m_write_write :  STD_LOGIC;
                signal sgdma_rx_m_write_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_csr_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sgdma_tx_csr_chipselect :  STD_LOGIC;
                signal sgdma_tx_csr_irq :  STD_LOGIC;
                signal sgdma_tx_csr_irq_from_sa :  STD_LOGIC;
                signal sgdma_tx_csr_read :  STD_LOGIC;
                signal sgdma_tx_csr_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_csr_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_csr_reset_n :  STD_LOGIC;
                signal sgdma_tx_csr_write :  STD_LOGIC;
                signal sgdma_tx_csr_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_read_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_latency_counter :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_read_readdatavalid :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_waitrequest :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_waitrequest :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_write :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_m_read_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_m_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_latency_counter :  STD_LOGIC;
                signal sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_read :  STD_LOGIC;
                signal sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1_shift_register :  STD_LOGIC;
                signal sgdma_tx_m_read_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_m_read_readdatavalid :  STD_LOGIC;
                signal sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_waitrequest :  STD_LOGIC;
                signal sgdma_tx_out_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_out_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sgdma_tx_out_endofpacket :  STD_LOGIC;
                signal sgdma_tx_out_error :  STD_LOGIC;
                signal sgdma_tx_out_ready :  STD_LOGIC;
                signal sgdma_tx_out_startofpacket :  STD_LOGIC;
                signal sgdma_tx_out_valid :  STD_LOGIC;
                signal sys_clk_timer_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sys_clk_timer_s1_chipselect :  STD_LOGIC;
                signal sys_clk_timer_s1_irq :  STD_LOGIC;
                signal sys_clk_timer_s1_irq_from_sa :  STD_LOGIC;
                signal sys_clk_timer_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sys_clk_timer_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sys_clk_timer_s1_reset_n :  STD_LOGIC;
                signal sys_clk_timer_s1_write_n :  STD_LOGIC;
                signal sys_clk_timer_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sysid_control_slave_address :  STD_LOGIC;
                signal sysid_control_slave_clock :  STD_LOGIC;
                signal sysid_control_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_reset_n :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal tse_ddr_clock_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal tse_ddr_clock_bridge_m1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tse_ddr_clock_bridge_m1_endofpacket :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_granted_sdram_s1 :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_latency_counter :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_read :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1 :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_ddr_clock_bridge_m1_readdatavalid :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_requests_sdram_s1 :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_reset_n :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_waitrequest :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_write :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_endofpacket :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_read :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_readdatavalid :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_reset_n :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_waitrequest :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_write :  STD_LOGIC;
                signal tse_ddr_clock_bridge_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_control_port_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal tse_mac_control_port_read :  STD_LOGIC;
                signal tse_mac_control_port_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_control_port_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_control_port_reset :  STD_LOGIC;
                signal tse_mac_control_port_waitrequest :  STD_LOGIC;
                signal tse_mac_control_port_waitrequest_from_sa :  STD_LOGIC;
                signal tse_mac_control_port_write :  STD_LOGIC;
                signal tse_mac_control_port_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_receive_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_receive_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tse_mac_receive_endofpacket :  STD_LOGIC;
                signal tse_mac_receive_error :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal tse_mac_receive_ready :  STD_LOGIC;
                signal tse_mac_receive_startofpacket :  STD_LOGIC;
                signal tse_mac_receive_valid :  STD_LOGIC;
                signal tse_mac_transmit_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_transmit_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tse_mac_transmit_endofpacket :  STD_LOGIC;
                signal tse_mac_transmit_error :  STD_LOGIC;
                signal tse_mac_transmit_ready :  STD_LOGIC;
                signal tse_mac_transmit_ready_from_sa :  STD_LOGIC;
                signal tse_mac_transmit_startofpacket :  STD_LOGIC;
                signal tse_mac_transmit_valid :  STD_LOGIC;

begin

  --the_cpuNios_jtag_debug_module, which is an e_instance
  the_cpuNios_jtag_debug_module : cpuNios_jtag_debug_module_arbitrator
    port map(
      cpuNios_data_master_granted_cpuNios_jtag_debug_module => cpuNios_data_master_granted_cpuNios_jtag_debug_module,
      cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module => cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module,
      cpuNios_data_master_read_data_valid_cpuNios_jtag_debug_module => cpuNios_data_master_read_data_valid_cpuNios_jtag_debug_module,
      cpuNios_data_master_requests_cpuNios_jtag_debug_module => cpuNios_data_master_requests_cpuNios_jtag_debug_module,
      cpuNios_instruction_master_granted_cpuNios_jtag_debug_module => cpuNios_instruction_master_granted_cpuNios_jtag_debug_module,
      cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module => cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module,
      cpuNios_instruction_master_read_data_valid_cpuNios_jtag_debug_module => cpuNios_instruction_master_read_data_valid_cpuNios_jtag_debug_module,
      cpuNios_instruction_master_requests_cpuNios_jtag_debug_module => cpuNios_instruction_master_requests_cpuNios_jtag_debug_module,
      cpuNios_jtag_debug_module_address => cpuNios_jtag_debug_module_address,
      cpuNios_jtag_debug_module_begintransfer => cpuNios_jtag_debug_module_begintransfer,
      cpuNios_jtag_debug_module_byteenable => cpuNios_jtag_debug_module_byteenable,
      cpuNios_jtag_debug_module_chipselect => cpuNios_jtag_debug_module_chipselect,
      cpuNios_jtag_debug_module_debugaccess => cpuNios_jtag_debug_module_debugaccess,
      cpuNios_jtag_debug_module_readdata_from_sa => cpuNios_jtag_debug_module_readdata_from_sa,
      cpuNios_jtag_debug_module_reset_n => cpuNios_jtag_debug_module_reset_n,
      cpuNios_jtag_debug_module_resetrequest_from_sa => cpuNios_jtag_debug_module_resetrequest_from_sa,
      cpuNios_jtag_debug_module_write => cpuNios_jtag_debug_module_write,
      cpuNios_jtag_debug_module_writedata => cpuNios_jtag_debug_module_writedata,
      d1_cpuNios_jtag_debug_module_end_xfer => d1_cpuNios_jtag_debug_module_end_xfer,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_byteenable => cpuNios_data_master_byteenable,
      cpuNios_data_master_debugaccess => cpuNios_data_master_debugaccess,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      cpuNios_instruction_master_address_to_slave => cpuNios_instruction_master_address_to_slave,
      cpuNios_instruction_master_read => cpuNios_instruction_master_read,
      cpuNios_jtag_debug_module_readdata => cpuNios_jtag_debug_module_readdata,
      cpuNios_jtag_debug_module_resetrequest => cpuNios_jtag_debug_module_resetrequest,
      reset_n => clk100MHz_reset_n
    );


  --the_cpuNios_data_master, which is an e_instance
  the_cpuNios_data_master : cpuNios_data_master_arbitrator
    port map(
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_irq => cpuNios_data_master_irq,
      cpuNios_data_master_readdata => cpuNios_data_master_readdata,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      clk => clk100MHz,
      clk100MHz => clk100MHz,
      clk100MHz_reset_n => clk100MHz_reset_n,
      cpuNios_data_master_address => cpuNios_data_master_address,
      cpuNios_data_master_granted_cpuNios_jtag_debug_module => cpuNios_data_master_granted_cpuNios_jtag_debug_module,
      cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 => cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1,
      cpuNios_data_master_granted_descriptor_memory_s1 => cpuNios_data_master_granted_descriptor_memory_s1,
      cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 => cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0,
      cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave => cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave,
      cpuNios_data_master_granted_lcd_i2c_en_s1 => cpuNios_data_master_granted_lcd_i2c_en_s1,
      cpuNios_data_master_granted_lcd_i2c_scl_s1 => cpuNios_data_master_granted_lcd_i2c_scl_s1,
      cpuNios_data_master_granted_lcd_i2c_sdat_s1 => cpuNios_data_master_granted_lcd_i2c_sdat_s1,
      cpuNios_data_master_granted_performance_counter_control_slave => cpuNios_data_master_granted_performance_counter_control_slave,
      cpuNios_data_master_granted_sgdma_rx_csr => cpuNios_data_master_granted_sgdma_rx_csr,
      cpuNios_data_master_granted_sgdma_tx_csr => cpuNios_data_master_granted_sgdma_tx_csr,
      cpuNios_data_master_granted_sys_clk_timer_s1 => cpuNios_data_master_granted_sys_clk_timer_s1,
      cpuNios_data_master_granted_sysid_control_slave => cpuNios_data_master_granted_sysid_control_slave,
      cpuNios_data_master_granted_tse_mac_control_port => cpuNios_data_master_granted_tse_mac_control_port,
      cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module => cpuNios_data_master_qualified_request_cpuNios_jtag_debug_module,
      cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 => cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1,
      cpuNios_data_master_qualified_request_descriptor_memory_s1 => cpuNios_data_master_qualified_request_descriptor_memory_s1,
      cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 => cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0,
      cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave => cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave,
      cpuNios_data_master_qualified_request_lcd_i2c_en_s1 => cpuNios_data_master_qualified_request_lcd_i2c_en_s1,
      cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 => cpuNios_data_master_qualified_request_lcd_i2c_scl_s1,
      cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 => cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1,
      cpuNios_data_master_qualified_request_performance_counter_control_slave => cpuNios_data_master_qualified_request_performance_counter_control_slave,
      cpuNios_data_master_qualified_request_sgdma_rx_csr => cpuNios_data_master_qualified_request_sgdma_rx_csr,
      cpuNios_data_master_qualified_request_sgdma_tx_csr => cpuNios_data_master_qualified_request_sgdma_tx_csr,
      cpuNios_data_master_qualified_request_sys_clk_timer_s1 => cpuNios_data_master_qualified_request_sys_clk_timer_s1,
      cpuNios_data_master_qualified_request_sysid_control_slave => cpuNios_data_master_qualified_request_sysid_control_slave,
      cpuNios_data_master_qualified_request_tse_mac_control_port => cpuNios_data_master_qualified_request_tse_mac_control_port,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_read_data_valid_cpuNios_jtag_debug_module => cpuNios_data_master_read_data_valid_cpuNios_jtag_debug_module,
      cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 => cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1,
      cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register => cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
      cpuNios_data_master_read_data_valid_descriptor_memory_s1 => cpuNios_data_master_read_data_valid_descriptor_memory_s1,
      cpuNios_data_master_read_data_valid_fft_pipeline_0_avalon_slave_0 => cpuNios_data_master_read_data_valid_fft_pipeline_0_avalon_slave_0,
      cpuNios_data_master_read_data_valid_jtag_uart_avalon_jtag_slave => cpuNios_data_master_read_data_valid_jtag_uart_avalon_jtag_slave,
      cpuNios_data_master_read_data_valid_lcd_i2c_en_s1 => cpuNios_data_master_read_data_valid_lcd_i2c_en_s1,
      cpuNios_data_master_read_data_valid_lcd_i2c_scl_s1 => cpuNios_data_master_read_data_valid_lcd_i2c_scl_s1,
      cpuNios_data_master_read_data_valid_lcd_i2c_sdat_s1 => cpuNios_data_master_read_data_valid_lcd_i2c_sdat_s1,
      cpuNios_data_master_read_data_valid_performance_counter_control_slave => cpuNios_data_master_read_data_valid_performance_counter_control_slave,
      cpuNios_data_master_read_data_valid_sgdma_rx_csr => cpuNios_data_master_read_data_valid_sgdma_rx_csr,
      cpuNios_data_master_read_data_valid_sgdma_tx_csr => cpuNios_data_master_read_data_valid_sgdma_tx_csr,
      cpuNios_data_master_read_data_valid_sys_clk_timer_s1 => cpuNios_data_master_read_data_valid_sys_clk_timer_s1,
      cpuNios_data_master_read_data_valid_sysid_control_slave => cpuNios_data_master_read_data_valid_sysid_control_slave,
      cpuNios_data_master_read_data_valid_tse_mac_control_port => cpuNios_data_master_read_data_valid_tse_mac_control_port,
      cpuNios_data_master_requests_cpuNios_jtag_debug_module => cpuNios_data_master_requests_cpuNios_jtag_debug_module,
      cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 => cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1,
      cpuNios_data_master_requests_descriptor_memory_s1 => cpuNios_data_master_requests_descriptor_memory_s1,
      cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 => cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0,
      cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave => cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave,
      cpuNios_data_master_requests_lcd_i2c_en_s1 => cpuNios_data_master_requests_lcd_i2c_en_s1,
      cpuNios_data_master_requests_lcd_i2c_scl_s1 => cpuNios_data_master_requests_lcd_i2c_scl_s1,
      cpuNios_data_master_requests_lcd_i2c_sdat_s1 => cpuNios_data_master_requests_lcd_i2c_sdat_s1,
      cpuNios_data_master_requests_performance_counter_control_slave => cpuNios_data_master_requests_performance_counter_control_slave,
      cpuNios_data_master_requests_sgdma_rx_csr => cpuNios_data_master_requests_sgdma_rx_csr,
      cpuNios_data_master_requests_sgdma_tx_csr => cpuNios_data_master_requests_sgdma_tx_csr,
      cpuNios_data_master_requests_sys_clk_timer_s1 => cpuNios_data_master_requests_sys_clk_timer_s1,
      cpuNios_data_master_requests_sysid_control_slave => cpuNios_data_master_requests_sysid_control_slave,
      cpuNios_data_master_requests_tse_mac_control_port => cpuNios_data_master_requests_tse_mac_control_port,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_jtag_debug_module_readdata_from_sa => cpuNios_jtag_debug_module_readdata_from_sa,
      cpu_ddr_clock_bridge_s1_readdata_from_sa => cpu_ddr_clock_bridge_s1_readdata_from_sa,
      cpu_ddr_clock_bridge_s1_waitrequest_from_sa => cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
      d1_cpuNios_jtag_debug_module_end_xfer => d1_cpuNios_jtag_debug_module_end_xfer,
      d1_cpu_ddr_clock_bridge_s1_end_xfer => d1_cpu_ddr_clock_bridge_s1_end_xfer,
      d1_descriptor_memory_s1_end_xfer => d1_descriptor_memory_s1_end_xfer,
      d1_fft_pipeline_0_avalon_slave_0_end_xfer => d1_fft_pipeline_0_avalon_slave_0_end_xfer,
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      d1_lcd_i2c_en_s1_end_xfer => d1_lcd_i2c_en_s1_end_xfer,
      d1_lcd_i2c_scl_s1_end_xfer => d1_lcd_i2c_scl_s1_end_xfer,
      d1_lcd_i2c_sdat_s1_end_xfer => d1_lcd_i2c_sdat_s1_end_xfer,
      d1_performance_counter_control_slave_end_xfer => d1_performance_counter_control_slave_end_xfer,
      d1_sgdma_rx_csr_end_xfer => d1_sgdma_rx_csr_end_xfer,
      d1_sgdma_tx_csr_end_xfer => d1_sgdma_tx_csr_end_xfer,
      d1_sys_clk_timer_s1_end_xfer => d1_sys_clk_timer_s1_end_xfer,
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      d1_tse_mac_control_port_end_xfer => d1_tse_mac_control_port_end_xfer,
      descriptor_memory_s1_readdata_from_sa => descriptor_memory_s1_readdata_from_sa,
      fft_pipeline_0_avalon_slave_0_readdata_from_sa => fft_pipeline_0_avalon_slave_0_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      lcd_i2c_en_s1_readdata_from_sa => lcd_i2c_en_s1_readdata_from_sa,
      lcd_i2c_scl_s1_readdata_from_sa => lcd_i2c_scl_s1_readdata_from_sa,
      lcd_i2c_sdat_s1_readdata_from_sa => lcd_i2c_sdat_s1_readdata_from_sa,
      lcd_sgdma_csr_irq_from_sa => lcd_sgdma_csr_irq_from_sa,
      performance_counter_control_slave_readdata_from_sa => performance_counter_control_slave_readdata_from_sa,
      registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1 => registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1,
      registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave => registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave,
      reset_n => clk100MHz_reset_n,
      sgdma_rx_csr_irq_from_sa => sgdma_rx_csr_irq_from_sa,
      sgdma_rx_csr_readdata_from_sa => sgdma_rx_csr_readdata_from_sa,
      sgdma_tx_csr_irq_from_sa => sgdma_tx_csr_irq_from_sa,
      sgdma_tx_csr_readdata_from_sa => sgdma_tx_csr_readdata_from_sa,
      sys_clk_timer_s1_irq_from_sa => sys_clk_timer_s1_irq_from_sa,
      sys_clk_timer_s1_readdata_from_sa => sys_clk_timer_s1_readdata_from_sa,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa,
      tse_mac_control_port_readdata_from_sa => tse_mac_control_port_readdata_from_sa,
      tse_mac_control_port_waitrequest_from_sa => tse_mac_control_port_waitrequest_from_sa
    );


  --the_cpuNios_instruction_master, which is an e_instance
  the_cpuNios_instruction_master : cpuNios_instruction_master_arbitrator
    port map(
      cpuNios_instruction_master_address_to_slave => cpuNios_instruction_master_address_to_slave,
      cpuNios_instruction_master_readdata => cpuNios_instruction_master_readdata,
      cpuNios_instruction_master_waitrequest => cpuNios_instruction_master_waitrequest,
      clk => clk100MHz,
      cpuNios_instruction_master_address => cpuNios_instruction_master_address,
      cpuNios_instruction_master_granted_cpuNios_jtag_debug_module => cpuNios_instruction_master_granted_cpuNios_jtag_debug_module,
      cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 => cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1,
      cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module => cpuNios_instruction_master_qualified_request_cpuNios_jtag_debug_module,
      cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 => cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1,
      cpuNios_instruction_master_read => cpuNios_instruction_master_read,
      cpuNios_instruction_master_read_data_valid_cpuNios_jtag_debug_module => cpuNios_instruction_master_read_data_valid_cpuNios_jtag_debug_module,
      cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 => cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1,
      cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register => cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
      cpuNios_instruction_master_requests_cpuNios_jtag_debug_module => cpuNios_instruction_master_requests_cpuNios_jtag_debug_module,
      cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 => cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1,
      cpuNios_jtag_debug_module_readdata_from_sa => cpuNios_jtag_debug_module_readdata_from_sa,
      cpu_ddr_clock_bridge_s1_readdata_from_sa => cpu_ddr_clock_bridge_s1_readdata_from_sa,
      cpu_ddr_clock_bridge_s1_waitrequest_from_sa => cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
      d1_cpuNios_jtag_debug_module_end_xfer => d1_cpuNios_jtag_debug_module_end_xfer,
      d1_cpu_ddr_clock_bridge_s1_end_xfer => d1_cpu_ddr_clock_bridge_s1_end_xfer,
      reset_n => clk100MHz_reset_n
    );


  --the_cpuNios, which is an e_ptf_instance
  the_cpuNios : cpuNios
    port map(
      d_address => cpuNios_data_master_address,
      d_byteenable => cpuNios_data_master_byteenable,
      d_read => cpuNios_data_master_read,
      d_write => cpuNios_data_master_write,
      d_writedata => cpuNios_data_master_writedata,
      i_address => cpuNios_instruction_master_address,
      i_read => cpuNios_instruction_master_read,
      jtag_debug_module_debugaccess_to_roms => cpuNios_data_master_debugaccess,
      jtag_debug_module_readdata => cpuNios_jtag_debug_module_readdata,
      jtag_debug_module_resetrequest => cpuNios_jtag_debug_module_resetrequest,
      clk => clk100MHz,
      d_irq => cpuNios_data_master_irq,
      d_readdata => cpuNios_data_master_readdata,
      d_waitrequest => cpuNios_data_master_waitrequest,
      i_readdata => cpuNios_instruction_master_readdata,
      i_waitrequest => cpuNios_instruction_master_waitrequest,
      jtag_debug_module_address => cpuNios_jtag_debug_module_address,
      jtag_debug_module_begintransfer => cpuNios_jtag_debug_module_begintransfer,
      jtag_debug_module_byteenable => cpuNios_jtag_debug_module_byteenable,
      jtag_debug_module_debugaccess => cpuNios_jtag_debug_module_debugaccess,
      jtag_debug_module_select => cpuNios_jtag_debug_module_chipselect,
      jtag_debug_module_write => cpuNios_jtag_debug_module_write,
      jtag_debug_module_writedata => cpuNios_jtag_debug_module_writedata,
      reset_n => cpuNios_jtag_debug_module_reset_n
    );


  --the_cpu_ddr_clock_bridge_s1, which is an e_instance
  the_cpu_ddr_clock_bridge_s1 : cpu_ddr_clock_bridge_s1_arbitrator
    port map(
      cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1 => cpuNios_data_master_granted_cpu_ddr_clock_bridge_s1,
      cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1 => cpuNios_data_master_qualified_request_cpu_ddr_clock_bridge_s1,
      cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 => cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1,
      cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register => cpuNios_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
      cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1 => cpuNios_data_master_requests_cpu_ddr_clock_bridge_s1,
      cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1 => cpuNios_instruction_master_granted_cpu_ddr_clock_bridge_s1,
      cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 => cpuNios_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1,
      cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 => cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1,
      cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register => cpuNios_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
      cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1 => cpuNios_instruction_master_requests_cpu_ddr_clock_bridge_s1,
      cpu_ddr_clock_bridge_s1_address => cpu_ddr_clock_bridge_s1_address,
      cpu_ddr_clock_bridge_s1_byteenable => cpu_ddr_clock_bridge_s1_byteenable,
      cpu_ddr_clock_bridge_s1_endofpacket_from_sa => cpu_ddr_clock_bridge_s1_endofpacket_from_sa,
      cpu_ddr_clock_bridge_s1_nativeaddress => cpu_ddr_clock_bridge_s1_nativeaddress,
      cpu_ddr_clock_bridge_s1_read => cpu_ddr_clock_bridge_s1_read,
      cpu_ddr_clock_bridge_s1_readdata_from_sa => cpu_ddr_clock_bridge_s1_readdata_from_sa,
      cpu_ddr_clock_bridge_s1_reset_n => cpu_ddr_clock_bridge_s1_reset_n,
      cpu_ddr_clock_bridge_s1_waitrequest_from_sa => cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
      cpu_ddr_clock_bridge_s1_write => cpu_ddr_clock_bridge_s1_write,
      cpu_ddr_clock_bridge_s1_writedata => cpu_ddr_clock_bridge_s1_writedata,
      d1_cpu_ddr_clock_bridge_s1_end_xfer => d1_cpu_ddr_clock_bridge_s1_end_xfer,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_byteenable => cpuNios_data_master_byteenable,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      cpuNios_instruction_master_address_to_slave => cpuNios_instruction_master_address_to_slave,
      cpuNios_instruction_master_read => cpuNios_instruction_master_read,
      cpu_ddr_clock_bridge_s1_endofpacket => cpu_ddr_clock_bridge_s1_endofpacket,
      cpu_ddr_clock_bridge_s1_readdata => cpu_ddr_clock_bridge_s1_readdata,
      cpu_ddr_clock_bridge_s1_readdatavalid => cpu_ddr_clock_bridge_s1_readdatavalid,
      cpu_ddr_clock_bridge_s1_waitrequest => cpu_ddr_clock_bridge_s1_waitrequest,
      reset_n => clk100MHz_reset_n
    );


  --the_cpu_ddr_clock_bridge_m1, which is an e_instance
  the_cpu_ddr_clock_bridge_m1 : cpu_ddr_clock_bridge_m1_arbitrator
    port map(
      cpu_ddr_clock_bridge_m1_address_to_slave => cpu_ddr_clock_bridge_m1_address_to_slave,
      cpu_ddr_clock_bridge_m1_latency_counter => cpu_ddr_clock_bridge_m1_latency_counter,
      cpu_ddr_clock_bridge_m1_readdata => cpu_ddr_clock_bridge_m1_readdata,
      cpu_ddr_clock_bridge_m1_readdatavalid => cpu_ddr_clock_bridge_m1_readdatavalid,
      cpu_ddr_clock_bridge_m1_reset_n => cpu_ddr_clock_bridge_m1_reset_n,
      cpu_ddr_clock_bridge_m1_waitrequest => cpu_ddr_clock_bridge_m1_waitrequest,
      clk => internal_sdram_phy_clk_out,
      cpu_ddr_clock_bridge_m1_address => cpu_ddr_clock_bridge_m1_address,
      cpu_ddr_clock_bridge_m1_byteenable => cpu_ddr_clock_bridge_m1_byteenable,
      cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr => cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr,
      cpu_ddr_clock_bridge_m1_granted_sdram_s1 => cpu_ddr_clock_bridge_m1_granted_sdram_s1,
      cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr => cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr,
      cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 => cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1,
      cpu_ddr_clock_bridge_m1_read => cpu_ddr_clock_bridge_m1_read,
      cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr => cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr,
      cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1 => cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1,
      cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register => cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register,
      cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr => cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr,
      cpu_ddr_clock_bridge_m1_requests_sdram_s1 => cpu_ddr_clock_bridge_m1_requests_sdram_s1,
      cpu_ddr_clock_bridge_m1_write => cpu_ddr_clock_bridge_m1_write,
      cpu_ddr_clock_bridge_m1_writedata => cpu_ddr_clock_bridge_m1_writedata,
      d1_lcd_sgdma_csr_end_xfer => d1_lcd_sgdma_csr_end_xfer,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      lcd_sgdma_csr_readdata_from_sa => lcd_sgdma_csr_readdata_from_sa,
      reset_n => sdram_phy_clk_out_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_n_from_sa => sdram_s1_waitrequest_n_from_sa
    );


  --the_cpu_ddr_clock_bridge, which is an e_ptf_instance
  the_cpu_ddr_clock_bridge : cpu_ddr_clock_bridge
    port map(
      master_address => cpu_ddr_clock_bridge_m1_address,
      master_byteenable => cpu_ddr_clock_bridge_m1_byteenable,
      master_nativeaddress => cpu_ddr_clock_bridge_m1_nativeaddress,
      master_read => cpu_ddr_clock_bridge_m1_read,
      master_write => cpu_ddr_clock_bridge_m1_write,
      master_writedata => cpu_ddr_clock_bridge_m1_writedata,
      slave_endofpacket => cpu_ddr_clock_bridge_s1_endofpacket,
      slave_readdata => cpu_ddr_clock_bridge_s1_readdata,
      slave_readdatavalid => cpu_ddr_clock_bridge_s1_readdatavalid,
      slave_waitrequest => cpu_ddr_clock_bridge_s1_waitrequest,
      master_clk => internal_sdram_phy_clk_out,
      master_endofpacket => cpu_ddr_clock_bridge_m1_endofpacket,
      master_readdata => cpu_ddr_clock_bridge_m1_readdata,
      master_readdatavalid => cpu_ddr_clock_bridge_m1_readdatavalid,
      master_reset_n => cpu_ddr_clock_bridge_m1_reset_n,
      master_waitrequest => cpu_ddr_clock_bridge_m1_waitrequest,
      slave_address => cpu_ddr_clock_bridge_s1_address,
      slave_byteenable => cpu_ddr_clock_bridge_s1_byteenable,
      slave_clk => clk100MHz,
      slave_nativeaddress => cpu_ddr_clock_bridge_s1_nativeaddress,
      slave_read => cpu_ddr_clock_bridge_s1_read,
      slave_reset_n => cpu_ddr_clock_bridge_s1_reset_n,
      slave_write => cpu_ddr_clock_bridge_s1_write,
      slave_writedata => cpu_ddr_clock_bridge_s1_writedata
    );


  --the_descriptor_memory_s1, which is an e_instance
  the_descriptor_memory_s1 : descriptor_memory_s1_arbitrator
    port map(
      cpuNios_data_master_granted_descriptor_memory_s1 => cpuNios_data_master_granted_descriptor_memory_s1,
      cpuNios_data_master_qualified_request_descriptor_memory_s1 => cpuNios_data_master_qualified_request_descriptor_memory_s1,
      cpuNios_data_master_read_data_valid_descriptor_memory_s1 => cpuNios_data_master_read_data_valid_descriptor_memory_s1,
      cpuNios_data_master_requests_descriptor_memory_s1 => cpuNios_data_master_requests_descriptor_memory_s1,
      d1_descriptor_memory_s1_end_xfer => d1_descriptor_memory_s1_end_xfer,
      descriptor_memory_s1_address => descriptor_memory_s1_address,
      descriptor_memory_s1_byteenable => descriptor_memory_s1_byteenable,
      descriptor_memory_s1_chipselect => descriptor_memory_s1_chipselect,
      descriptor_memory_s1_clken => descriptor_memory_s1_clken,
      descriptor_memory_s1_readdata_from_sa => descriptor_memory_s1_readdata_from_sa,
      descriptor_memory_s1_reset => descriptor_memory_s1_reset,
      descriptor_memory_s1_write => descriptor_memory_s1_write,
      descriptor_memory_s1_writedata => descriptor_memory_s1_writedata,
      descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1 => descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1,
      descriptor_offset_bridge_m1_granted_descriptor_memory_s1 => descriptor_offset_bridge_m1_granted_descriptor_memory_s1,
      descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 => descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1,
      descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1 => descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1,
      descriptor_offset_bridge_m1_requests_descriptor_memory_s1 => descriptor_offset_bridge_m1_requests_descriptor_memory_s1,
      registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1 => registered_cpuNios_data_master_read_data_valid_descriptor_memory_s1,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_byteenable => cpuNios_data_master_byteenable,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      descriptor_memory_s1_readdata => descriptor_memory_s1_readdata,
      descriptor_offset_bridge_m1_address_to_slave => descriptor_offset_bridge_m1_address_to_slave,
      descriptor_offset_bridge_m1_burstcount => descriptor_offset_bridge_m1_burstcount,
      descriptor_offset_bridge_m1_byteenable => descriptor_offset_bridge_m1_byteenable,
      descriptor_offset_bridge_m1_chipselect => descriptor_offset_bridge_m1_chipselect,
      descriptor_offset_bridge_m1_dbs_address => descriptor_offset_bridge_m1_dbs_address,
      descriptor_offset_bridge_m1_dbs_write_32 => descriptor_offset_bridge_m1_dbs_write_32,
      descriptor_offset_bridge_m1_latency_counter => descriptor_offset_bridge_m1_latency_counter,
      descriptor_offset_bridge_m1_read => descriptor_offset_bridge_m1_read,
      descriptor_offset_bridge_m1_write => descriptor_offset_bridge_m1_write,
      reset_n => clk100MHz_reset_n
    );


  --the_descriptor_memory, which is an e_ptf_instance
  the_descriptor_memory : descriptor_memory
    port map(
      readdata => descriptor_memory_s1_readdata,
      address => descriptor_memory_s1_address,
      byteenable => descriptor_memory_s1_byteenable,
      chipselect => descriptor_memory_s1_chipselect,
      clk => clk100MHz,
      clken => descriptor_memory_s1_clken,
      reset => descriptor_memory_s1_reset,
      write => descriptor_memory_s1_write,
      writedata => descriptor_memory_s1_writedata
    );


  --the_descriptor_offset_bridge_s1, which is an e_instance
  the_descriptor_offset_bridge_s1 : descriptor_offset_bridge_s1_arbitrator
    port map(
      d1_descriptor_offset_bridge_s1_end_xfer => d1_descriptor_offset_bridge_s1_end_xfer,
      descriptor_offset_bridge_s1_address => descriptor_offset_bridge_s1_address,
      descriptor_offset_bridge_s1_arbiterlock => descriptor_offset_bridge_s1_arbiterlock,
      descriptor_offset_bridge_s1_arbiterlock2 => descriptor_offset_bridge_s1_arbiterlock2,
      descriptor_offset_bridge_s1_burstcount => descriptor_offset_bridge_s1_burstcount,
      descriptor_offset_bridge_s1_byteenable => descriptor_offset_bridge_s1_byteenable,
      descriptor_offset_bridge_s1_chipselect => descriptor_offset_bridge_s1_chipselect,
      descriptor_offset_bridge_s1_debugaccess => descriptor_offset_bridge_s1_debugaccess,
      descriptor_offset_bridge_s1_endofpacket_from_sa => descriptor_offset_bridge_s1_endofpacket_from_sa,
      descriptor_offset_bridge_s1_nativeaddress => descriptor_offset_bridge_s1_nativeaddress,
      descriptor_offset_bridge_s1_read => descriptor_offset_bridge_s1_read,
      descriptor_offset_bridge_s1_readdata_from_sa => descriptor_offset_bridge_s1_readdata_from_sa,
      descriptor_offset_bridge_s1_reset_n => descriptor_offset_bridge_s1_reset_n,
      descriptor_offset_bridge_s1_waitrequest_from_sa => descriptor_offset_bridge_s1_waitrequest_from_sa,
      descriptor_offset_bridge_s1_write => descriptor_offset_bridge_s1_write,
      descriptor_offset_bridge_s1_writedata => descriptor_offset_bridge_s1_writedata,
      sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register => sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register,
      sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register => sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register,
      sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1,
      clk => clk100MHz,
      descriptor_offset_bridge_s1_endofpacket => descriptor_offset_bridge_s1_endofpacket,
      descriptor_offset_bridge_s1_readdata => descriptor_offset_bridge_s1_readdata,
      descriptor_offset_bridge_s1_readdatavalid => descriptor_offset_bridge_s1_readdatavalid,
      descriptor_offset_bridge_s1_waitrequest => descriptor_offset_bridge_s1_waitrequest,
      reset_n => clk100MHz_reset_n,
      sgdma_rx_descriptor_read_address_to_slave => sgdma_rx_descriptor_read_address_to_slave,
      sgdma_rx_descriptor_read_latency_counter => sgdma_rx_descriptor_read_latency_counter,
      sgdma_rx_descriptor_read_read => sgdma_rx_descriptor_read_read,
      sgdma_rx_descriptor_write_address_to_slave => sgdma_rx_descriptor_write_address_to_slave,
      sgdma_rx_descriptor_write_write => sgdma_rx_descriptor_write_write,
      sgdma_rx_descriptor_write_writedata => sgdma_rx_descriptor_write_writedata,
      sgdma_tx_descriptor_read_address_to_slave => sgdma_tx_descriptor_read_address_to_slave,
      sgdma_tx_descriptor_read_latency_counter => sgdma_tx_descriptor_read_latency_counter,
      sgdma_tx_descriptor_read_read => sgdma_tx_descriptor_read_read,
      sgdma_tx_descriptor_write_address_to_slave => sgdma_tx_descriptor_write_address_to_slave,
      sgdma_tx_descriptor_write_write => sgdma_tx_descriptor_write_write,
      sgdma_tx_descriptor_write_writedata => sgdma_tx_descriptor_write_writedata
    );


  --the_descriptor_offset_bridge_m1, which is an e_instance
  the_descriptor_offset_bridge_m1 : descriptor_offset_bridge_m1_arbitrator
    port map(
      descriptor_offset_bridge_m1_address_to_slave => descriptor_offset_bridge_m1_address_to_slave,
      descriptor_offset_bridge_m1_dbs_address => descriptor_offset_bridge_m1_dbs_address,
      descriptor_offset_bridge_m1_dbs_write_32 => descriptor_offset_bridge_m1_dbs_write_32,
      descriptor_offset_bridge_m1_latency_counter => descriptor_offset_bridge_m1_latency_counter,
      descriptor_offset_bridge_m1_readdata => descriptor_offset_bridge_m1_readdata,
      descriptor_offset_bridge_m1_readdatavalid => descriptor_offset_bridge_m1_readdatavalid,
      descriptor_offset_bridge_m1_waitrequest => descriptor_offset_bridge_m1_waitrequest,
      clk => clk100MHz,
      d1_descriptor_memory_s1_end_xfer => d1_descriptor_memory_s1_end_xfer,
      descriptor_memory_s1_readdata_from_sa => descriptor_memory_s1_readdata_from_sa,
      descriptor_offset_bridge_m1_address => descriptor_offset_bridge_m1_address,
      descriptor_offset_bridge_m1_burstcount => descriptor_offset_bridge_m1_burstcount,
      descriptor_offset_bridge_m1_byteenable => descriptor_offset_bridge_m1_byteenable,
      descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1 => descriptor_offset_bridge_m1_byteenable_descriptor_memory_s1,
      descriptor_offset_bridge_m1_chipselect => descriptor_offset_bridge_m1_chipselect,
      descriptor_offset_bridge_m1_granted_descriptor_memory_s1 => descriptor_offset_bridge_m1_granted_descriptor_memory_s1,
      descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1 => descriptor_offset_bridge_m1_qualified_request_descriptor_memory_s1,
      descriptor_offset_bridge_m1_read => descriptor_offset_bridge_m1_read,
      descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1 => descriptor_offset_bridge_m1_read_data_valid_descriptor_memory_s1,
      descriptor_offset_bridge_m1_requests_descriptor_memory_s1 => descriptor_offset_bridge_m1_requests_descriptor_memory_s1,
      descriptor_offset_bridge_m1_write => descriptor_offset_bridge_m1_write,
      descriptor_offset_bridge_m1_writedata => descriptor_offset_bridge_m1_writedata,
      reset_n => clk100MHz_reset_n
    );


  --the_descriptor_offset_bridge, which is an e_ptf_instance
  the_descriptor_offset_bridge : descriptor_offset_bridge
    port map(
      m1_address => descriptor_offset_bridge_m1_address,
      m1_burstcount => descriptor_offset_bridge_m1_burstcount,
      m1_byteenable => descriptor_offset_bridge_m1_byteenable,
      m1_chipselect => descriptor_offset_bridge_m1_chipselect,
      m1_debugaccess => descriptor_offset_bridge_m1_debugaccess,
      m1_read => descriptor_offset_bridge_m1_read,
      m1_write => descriptor_offset_bridge_m1_write,
      m1_writedata => descriptor_offset_bridge_m1_writedata,
      s1_endofpacket => descriptor_offset_bridge_s1_endofpacket,
      s1_readdata => descriptor_offset_bridge_s1_readdata,
      s1_readdatavalid => descriptor_offset_bridge_s1_readdatavalid,
      s1_waitrequest => descriptor_offset_bridge_s1_waitrequest,
      clk => clk100MHz,
      m1_endofpacket => descriptor_offset_bridge_m1_endofpacket,
      m1_readdata => descriptor_offset_bridge_m1_readdata,
      m1_readdatavalid => descriptor_offset_bridge_m1_readdatavalid,
      m1_waitrequest => descriptor_offset_bridge_m1_waitrequest,
      reset_n => descriptor_offset_bridge_s1_reset_n,
      s1_address => descriptor_offset_bridge_s1_address,
      s1_arbiterlock => descriptor_offset_bridge_s1_arbiterlock,
      s1_arbiterlock2 => descriptor_offset_bridge_s1_arbiterlock2,
      s1_burstcount => descriptor_offset_bridge_s1_burstcount,
      s1_byteenable => descriptor_offset_bridge_s1_byteenable,
      s1_chipselect => descriptor_offset_bridge_s1_chipselect,
      s1_debugaccess => descriptor_offset_bridge_s1_debugaccess,
      s1_nativeaddress => descriptor_offset_bridge_s1_nativeaddress,
      s1_read => descriptor_offset_bridge_s1_read,
      s1_write => descriptor_offset_bridge_s1_write,
      s1_writedata => descriptor_offset_bridge_s1_writedata
    );


  --the_fft_pipeline_0_avalon_slave_0, which is an e_instance
  the_fft_pipeline_0_avalon_slave_0 : fft_pipeline_0_avalon_slave_0_arbitrator
    port map(
      cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0 => cpuNios_data_master_granted_fft_pipeline_0_avalon_slave_0,
      cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0 => cpuNios_data_master_qualified_request_fft_pipeline_0_avalon_slave_0,
      cpuNios_data_master_read_data_valid_fft_pipeline_0_avalon_slave_0 => cpuNios_data_master_read_data_valid_fft_pipeline_0_avalon_slave_0,
      cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0 => cpuNios_data_master_requests_fft_pipeline_0_avalon_slave_0,
      d1_fft_pipeline_0_avalon_slave_0_end_xfer => d1_fft_pipeline_0_avalon_slave_0_end_xfer,
      fft_pipeline_0_avalon_slave_0_address => fft_pipeline_0_avalon_slave_0_address,
      fft_pipeline_0_avalon_slave_0_chipselect => fft_pipeline_0_avalon_slave_0_chipselect,
      fft_pipeline_0_avalon_slave_0_readdata_from_sa => fft_pipeline_0_avalon_slave_0_readdata_from_sa,
      fft_pipeline_0_avalon_slave_0_reset => fft_pipeline_0_avalon_slave_0_reset,
      fft_pipeline_0_avalon_slave_0_write => fft_pipeline_0_avalon_slave_0_write,
      fft_pipeline_0_avalon_slave_0_writedata => fft_pipeline_0_avalon_slave_0_writedata,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      fft_pipeline_0_avalon_slave_0_readdata => fft_pipeline_0_avalon_slave_0_readdata,
      reset_n => clk100MHz_reset_n
    );


  --the_fft_pipeline_0, which is an e_ptf_instance
  the_fft_pipeline_0 : fft_pipeline_0
    port map(
      counter => internal_counter_from_the_fft_pipeline_0,
      rd_data => fft_pipeline_0_avalon_slave_0_readdata,
      tx_out => internal_tx_out_from_the_fft_pipeline_0,
      addr => fft_pipeline_0_avalon_slave_0_address,
      clk => clk100MHz,
      clr_n => fft_pipeline_0_avalon_slave_0_reset,
      cs => fft_pipeline_0_avalon_slave_0_chipselect,
      rx_in => rx_in_to_the_fft_pipeline_0,
      wr => fft_pipeline_0_avalon_slave_0_write,
      wr_data => fft_pipeline_0_avalon_slave_0_writedata
    );


  --the_jtag_uart_avalon_jtag_slave, which is an e_instance
  the_jtag_uart_avalon_jtag_slave : jtag_uart_avalon_jtag_slave_arbitrator
    port map(
      cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave => cpuNios_data_master_granted_jtag_uart_avalon_jtag_slave,
      cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave => cpuNios_data_master_qualified_request_jtag_uart_avalon_jtag_slave,
      cpuNios_data_master_read_data_valid_jtag_uart_avalon_jtag_slave => cpuNios_data_master_read_data_valid_jtag_uart_avalon_jtag_slave,
      cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave => cpuNios_data_master_requests_jtag_uart_avalon_jtag_slave,
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      jtag_uart_avalon_jtag_slave_address => jtag_uart_avalon_jtag_slave_address,
      jtag_uart_avalon_jtag_slave_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      jtag_uart_avalon_jtag_slave_dataavailable_from_sa => jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      jtag_uart_avalon_jtag_slave_read_n => jtag_uart_avalon_jtag_slave_read_n,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_readyfordata_from_sa => jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
      jtag_uart_avalon_jtag_slave_reset_n => jtag_uart_avalon_jtag_slave_reset_n,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      jtag_uart_avalon_jtag_slave_write_n => jtag_uart_avalon_jtag_slave_write_n,
      jtag_uart_avalon_jtag_slave_writedata => jtag_uart_avalon_jtag_slave_writedata,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      jtag_uart_avalon_jtag_slave_dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      jtag_uart_avalon_jtag_slave_irq => jtag_uart_avalon_jtag_slave_irq,
      jtag_uart_avalon_jtag_slave_readdata => jtag_uart_avalon_jtag_slave_readdata,
      jtag_uart_avalon_jtag_slave_readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      jtag_uart_avalon_jtag_slave_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      reset_n => clk100MHz_reset_n
    );


  --the_jtag_uart, which is an e_ptf_instance
  the_jtag_uart : jtag_uart
    port map(
      av_irq => jtag_uart_avalon_jtag_slave_irq,
      av_readdata => jtag_uart_avalon_jtag_slave_readdata,
      av_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      av_address => jtag_uart_avalon_jtag_slave_address,
      av_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      av_read_n => jtag_uart_avalon_jtag_slave_read_n,
      av_write_n => jtag_uart_avalon_jtag_slave_write_n,
      av_writedata => jtag_uart_avalon_jtag_slave_writedata,
      clk => clk100MHz,
      rst_n => jtag_uart_avalon_jtag_slave_reset_n
    );


  --the_lcd_24_to_8_bits_dfa_in, which is an e_instance
  the_lcd_24_to_8_bits_dfa_in : lcd_24_to_8_bits_dfa_in_arbitrator
    port map(
      lcd_24_to_8_bits_dfa_in_data => lcd_24_to_8_bits_dfa_in_data,
      lcd_24_to_8_bits_dfa_in_empty => lcd_24_to_8_bits_dfa_in_empty,
      lcd_24_to_8_bits_dfa_in_endofpacket => lcd_24_to_8_bits_dfa_in_endofpacket,
      lcd_24_to_8_bits_dfa_in_ready_from_sa => lcd_24_to_8_bits_dfa_in_ready_from_sa,
      lcd_24_to_8_bits_dfa_in_reset_n => lcd_24_to_8_bits_dfa_in_reset_n,
      lcd_24_to_8_bits_dfa_in_startofpacket => lcd_24_to_8_bits_dfa_in_startofpacket,
      lcd_24_to_8_bits_dfa_in_valid => lcd_24_to_8_bits_dfa_in_valid,
      clk => clk100MHz,
      lcd_24_to_8_bits_dfa_in_ready => lcd_24_to_8_bits_dfa_in_ready,
      lcd_pixel_converter_out_data => lcd_pixel_converter_out_data,
      lcd_pixel_converter_out_empty => lcd_pixel_converter_out_empty,
      lcd_pixel_converter_out_endofpacket => lcd_pixel_converter_out_endofpacket,
      lcd_pixel_converter_out_startofpacket => lcd_pixel_converter_out_startofpacket,
      lcd_pixel_converter_out_valid => lcd_pixel_converter_out_valid,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_24_to_8_bits_dfa_out, which is an e_instance
  the_lcd_24_to_8_bits_dfa_out : lcd_24_to_8_bits_dfa_out_arbitrator
    port map(
      lcd_24_to_8_bits_dfa_out_ready => lcd_24_to_8_bits_dfa_out_ready,
      clk => clk100MHz,
      lcd_24_to_8_bits_dfa_out_data => lcd_24_to_8_bits_dfa_out_data,
      lcd_24_to_8_bits_dfa_out_empty => lcd_24_to_8_bits_dfa_out_empty,
      lcd_24_to_8_bits_dfa_out_endofpacket => lcd_24_to_8_bits_dfa_out_endofpacket,
      lcd_24_to_8_bits_dfa_out_startofpacket => lcd_24_to_8_bits_dfa_out_startofpacket,
      lcd_24_to_8_bits_dfa_out_valid => lcd_24_to_8_bits_dfa_out_valid,
      lcd_sync_generator_in_ready_from_sa => lcd_sync_generator_in_ready_from_sa,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_24_to_8_bits_dfa, which is an e_ptf_instance
  the_lcd_24_to_8_bits_dfa : lcd_24_to_8_bits_dfa
    port map(
      in_ready => lcd_24_to_8_bits_dfa_in_ready,
      out_data => lcd_24_to_8_bits_dfa_out_data,
      out_empty => lcd_24_to_8_bits_dfa_out_empty,
      out_endofpacket => lcd_24_to_8_bits_dfa_out_endofpacket,
      out_startofpacket => lcd_24_to_8_bits_dfa_out_startofpacket,
      out_valid => lcd_24_to_8_bits_dfa_out_valid,
      clk => clk100MHz,
      in_data => lcd_24_to_8_bits_dfa_in_data,
      in_empty => lcd_24_to_8_bits_dfa_in_empty,
      in_endofpacket => lcd_24_to_8_bits_dfa_in_endofpacket,
      in_startofpacket => lcd_24_to_8_bits_dfa_in_startofpacket,
      in_valid => lcd_24_to_8_bits_dfa_in_valid,
      out_ready => lcd_24_to_8_bits_dfa_out_ready,
      reset_n => lcd_24_to_8_bits_dfa_in_reset_n
    );


  --the_lcd_64_to_32_bits_dfa_in, which is an e_instance
  the_lcd_64_to_32_bits_dfa_in : lcd_64_to_32_bits_dfa_in_arbitrator
    port map(
      lcd_64_to_32_bits_dfa_in_data => lcd_64_to_32_bits_dfa_in_data,
      lcd_64_to_32_bits_dfa_in_empty => lcd_64_to_32_bits_dfa_in_empty,
      lcd_64_to_32_bits_dfa_in_endofpacket => lcd_64_to_32_bits_dfa_in_endofpacket,
      lcd_64_to_32_bits_dfa_in_ready_from_sa => lcd_64_to_32_bits_dfa_in_ready_from_sa,
      lcd_64_to_32_bits_dfa_in_reset_n => lcd_64_to_32_bits_dfa_in_reset_n,
      lcd_64_to_32_bits_dfa_in_startofpacket => lcd_64_to_32_bits_dfa_in_startofpacket,
      lcd_64_to_32_bits_dfa_in_valid => lcd_64_to_32_bits_dfa_in_valid,
      clk => clk100MHz,
      lcd_64_to_32_bits_dfa_in_ready => lcd_64_to_32_bits_dfa_in_ready,
      lcd_ta_fifo_to_dfa_out_data => lcd_ta_fifo_to_dfa_out_data,
      lcd_ta_fifo_to_dfa_out_empty => lcd_ta_fifo_to_dfa_out_empty,
      lcd_ta_fifo_to_dfa_out_endofpacket => lcd_ta_fifo_to_dfa_out_endofpacket,
      lcd_ta_fifo_to_dfa_out_startofpacket => lcd_ta_fifo_to_dfa_out_startofpacket,
      lcd_ta_fifo_to_dfa_out_valid => lcd_ta_fifo_to_dfa_out_valid,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_64_to_32_bits_dfa_out, which is an e_instance
  the_lcd_64_to_32_bits_dfa_out : lcd_64_to_32_bits_dfa_out_arbitrator
    port map(
      lcd_64_to_32_bits_dfa_out_ready => lcd_64_to_32_bits_dfa_out_ready,
      clk => clk100MHz,
      lcd_64_to_32_bits_dfa_out_data => lcd_64_to_32_bits_dfa_out_data,
      lcd_64_to_32_bits_dfa_out_empty => lcd_64_to_32_bits_dfa_out_empty,
      lcd_64_to_32_bits_dfa_out_endofpacket => lcd_64_to_32_bits_dfa_out_endofpacket,
      lcd_64_to_32_bits_dfa_out_startofpacket => lcd_64_to_32_bits_dfa_out_startofpacket,
      lcd_64_to_32_bits_dfa_out_valid => lcd_64_to_32_bits_dfa_out_valid,
      lcd_pixel_converter_in_ready_from_sa => lcd_pixel_converter_in_ready_from_sa,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_64_to_32_bits_dfa, which is an e_ptf_instance
  the_lcd_64_to_32_bits_dfa : lcd_64_to_32_bits_dfa
    port map(
      in_ready => lcd_64_to_32_bits_dfa_in_ready,
      out_data => lcd_64_to_32_bits_dfa_out_data,
      out_empty => lcd_64_to_32_bits_dfa_out_empty,
      out_endofpacket => lcd_64_to_32_bits_dfa_out_endofpacket,
      out_startofpacket => lcd_64_to_32_bits_dfa_out_startofpacket,
      out_valid => lcd_64_to_32_bits_dfa_out_valid,
      clk => clk100MHz,
      in_data => lcd_64_to_32_bits_dfa_in_data,
      in_empty => lcd_64_to_32_bits_dfa_in_empty,
      in_endofpacket => lcd_64_to_32_bits_dfa_in_endofpacket,
      in_startofpacket => lcd_64_to_32_bits_dfa_in_startofpacket,
      in_valid => lcd_64_to_32_bits_dfa_in_valid,
      out_ready => lcd_64_to_32_bits_dfa_out_ready,
      reset_n => lcd_64_to_32_bits_dfa_in_reset_n
    );


  --the_lcd_i2c_en_s1, which is an e_instance
  the_lcd_i2c_en_s1 : lcd_i2c_en_s1_arbitrator
    port map(
      cpuNios_data_master_granted_lcd_i2c_en_s1 => cpuNios_data_master_granted_lcd_i2c_en_s1,
      cpuNios_data_master_qualified_request_lcd_i2c_en_s1 => cpuNios_data_master_qualified_request_lcd_i2c_en_s1,
      cpuNios_data_master_read_data_valid_lcd_i2c_en_s1 => cpuNios_data_master_read_data_valid_lcd_i2c_en_s1,
      cpuNios_data_master_requests_lcd_i2c_en_s1 => cpuNios_data_master_requests_lcd_i2c_en_s1,
      d1_lcd_i2c_en_s1_end_xfer => d1_lcd_i2c_en_s1_end_xfer,
      lcd_i2c_en_s1_address => lcd_i2c_en_s1_address,
      lcd_i2c_en_s1_chipselect => lcd_i2c_en_s1_chipselect,
      lcd_i2c_en_s1_readdata_from_sa => lcd_i2c_en_s1_readdata_from_sa,
      lcd_i2c_en_s1_reset_n => lcd_i2c_en_s1_reset_n,
      lcd_i2c_en_s1_write_n => lcd_i2c_en_s1_write_n,
      lcd_i2c_en_s1_writedata => lcd_i2c_en_s1_writedata,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      lcd_i2c_en_s1_readdata => lcd_i2c_en_s1_readdata,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_i2c_en, which is an e_ptf_instance
  the_lcd_i2c_en : lcd_i2c_en
    port map(
      out_port => internal_out_port_from_the_lcd_i2c_en,
      readdata => lcd_i2c_en_s1_readdata,
      address => lcd_i2c_en_s1_address,
      chipselect => lcd_i2c_en_s1_chipselect,
      clk => clk100MHz,
      reset_n => lcd_i2c_en_s1_reset_n,
      write_n => lcd_i2c_en_s1_write_n,
      writedata => lcd_i2c_en_s1_writedata
    );


  --the_lcd_i2c_scl_s1, which is an e_instance
  the_lcd_i2c_scl_s1 : lcd_i2c_scl_s1_arbitrator
    port map(
      cpuNios_data_master_granted_lcd_i2c_scl_s1 => cpuNios_data_master_granted_lcd_i2c_scl_s1,
      cpuNios_data_master_qualified_request_lcd_i2c_scl_s1 => cpuNios_data_master_qualified_request_lcd_i2c_scl_s1,
      cpuNios_data_master_read_data_valid_lcd_i2c_scl_s1 => cpuNios_data_master_read_data_valid_lcd_i2c_scl_s1,
      cpuNios_data_master_requests_lcd_i2c_scl_s1 => cpuNios_data_master_requests_lcd_i2c_scl_s1,
      d1_lcd_i2c_scl_s1_end_xfer => d1_lcd_i2c_scl_s1_end_xfer,
      lcd_i2c_scl_s1_address => lcd_i2c_scl_s1_address,
      lcd_i2c_scl_s1_chipselect => lcd_i2c_scl_s1_chipselect,
      lcd_i2c_scl_s1_readdata_from_sa => lcd_i2c_scl_s1_readdata_from_sa,
      lcd_i2c_scl_s1_reset_n => lcd_i2c_scl_s1_reset_n,
      lcd_i2c_scl_s1_write_n => lcd_i2c_scl_s1_write_n,
      lcd_i2c_scl_s1_writedata => lcd_i2c_scl_s1_writedata,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      lcd_i2c_scl_s1_readdata => lcd_i2c_scl_s1_readdata,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_i2c_scl, which is an e_ptf_instance
  the_lcd_i2c_scl : lcd_i2c_scl
    port map(
      out_port => internal_out_port_from_the_lcd_i2c_scl,
      readdata => lcd_i2c_scl_s1_readdata,
      address => lcd_i2c_scl_s1_address,
      chipselect => lcd_i2c_scl_s1_chipselect,
      clk => clk100MHz,
      reset_n => lcd_i2c_scl_s1_reset_n,
      write_n => lcd_i2c_scl_s1_write_n,
      writedata => lcd_i2c_scl_s1_writedata
    );


  --the_lcd_i2c_sdat_s1, which is an e_instance
  the_lcd_i2c_sdat_s1 : lcd_i2c_sdat_s1_arbitrator
    port map(
      cpuNios_data_master_granted_lcd_i2c_sdat_s1 => cpuNios_data_master_granted_lcd_i2c_sdat_s1,
      cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1 => cpuNios_data_master_qualified_request_lcd_i2c_sdat_s1,
      cpuNios_data_master_read_data_valid_lcd_i2c_sdat_s1 => cpuNios_data_master_read_data_valid_lcd_i2c_sdat_s1,
      cpuNios_data_master_requests_lcd_i2c_sdat_s1 => cpuNios_data_master_requests_lcd_i2c_sdat_s1,
      d1_lcd_i2c_sdat_s1_end_xfer => d1_lcd_i2c_sdat_s1_end_xfer,
      lcd_i2c_sdat_s1_address => lcd_i2c_sdat_s1_address,
      lcd_i2c_sdat_s1_chipselect => lcd_i2c_sdat_s1_chipselect,
      lcd_i2c_sdat_s1_readdata_from_sa => lcd_i2c_sdat_s1_readdata_from_sa,
      lcd_i2c_sdat_s1_reset_n => lcd_i2c_sdat_s1_reset_n,
      lcd_i2c_sdat_s1_write_n => lcd_i2c_sdat_s1_write_n,
      lcd_i2c_sdat_s1_writedata => lcd_i2c_sdat_s1_writedata,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      lcd_i2c_sdat_s1_readdata => lcd_i2c_sdat_s1_readdata,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_i2c_sdat, which is an e_ptf_instance
  the_lcd_i2c_sdat : lcd_i2c_sdat
    port map(
      bidir_port => bidir_port_to_and_from_the_lcd_i2c_sdat,
      readdata => lcd_i2c_sdat_s1_readdata,
      address => lcd_i2c_sdat_s1_address,
      chipselect => lcd_i2c_sdat_s1_chipselect,
      clk => clk100MHz,
      reset_n => lcd_i2c_sdat_s1_reset_n,
      write_n => lcd_i2c_sdat_s1_write_n,
      writedata => lcd_i2c_sdat_s1_writedata
    );


  --the_lcd_pixel_converter_in, which is an e_instance
  the_lcd_pixel_converter_in : lcd_pixel_converter_in_arbitrator
    port map(
      lcd_pixel_converter_in_data => lcd_pixel_converter_in_data,
      lcd_pixel_converter_in_empty => lcd_pixel_converter_in_empty,
      lcd_pixel_converter_in_endofpacket => lcd_pixel_converter_in_endofpacket,
      lcd_pixel_converter_in_ready_from_sa => lcd_pixel_converter_in_ready_from_sa,
      lcd_pixel_converter_in_reset_n => lcd_pixel_converter_in_reset_n,
      lcd_pixel_converter_in_startofpacket => lcd_pixel_converter_in_startofpacket,
      lcd_pixel_converter_in_valid => lcd_pixel_converter_in_valid,
      clk => clk100MHz,
      lcd_64_to_32_bits_dfa_out_data => lcd_64_to_32_bits_dfa_out_data,
      lcd_64_to_32_bits_dfa_out_empty => lcd_64_to_32_bits_dfa_out_empty,
      lcd_64_to_32_bits_dfa_out_endofpacket => lcd_64_to_32_bits_dfa_out_endofpacket,
      lcd_64_to_32_bits_dfa_out_startofpacket => lcd_64_to_32_bits_dfa_out_startofpacket,
      lcd_64_to_32_bits_dfa_out_valid => lcd_64_to_32_bits_dfa_out_valid,
      lcd_pixel_converter_in_ready => lcd_pixel_converter_in_ready,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_pixel_converter_out, which is an e_instance
  the_lcd_pixel_converter_out : lcd_pixel_converter_out_arbitrator
    port map(
      lcd_pixel_converter_out_ready => lcd_pixel_converter_out_ready,
      clk => clk100MHz,
      lcd_24_to_8_bits_dfa_in_ready_from_sa => lcd_24_to_8_bits_dfa_in_ready_from_sa,
      lcd_pixel_converter_out_data => lcd_pixel_converter_out_data,
      lcd_pixel_converter_out_empty => lcd_pixel_converter_out_empty,
      lcd_pixel_converter_out_endofpacket => lcd_pixel_converter_out_endofpacket,
      lcd_pixel_converter_out_startofpacket => lcd_pixel_converter_out_startofpacket,
      lcd_pixel_converter_out_valid => lcd_pixel_converter_out_valid,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_pixel_converter, which is an e_ptf_instance
  the_lcd_pixel_converter : lcd_pixel_converter
    port map(
      data_out => lcd_pixel_converter_out_data,
      empty_out => lcd_pixel_converter_out_empty,
      eop_out => lcd_pixel_converter_out_endofpacket,
      ready_out => lcd_pixel_converter_in_ready,
      sop_out => lcd_pixel_converter_out_startofpacket,
      valid_out => lcd_pixel_converter_out_valid,
      clk => clk100MHz,
      data_in => lcd_pixel_converter_in_data,
      empty_in => lcd_pixel_converter_in_empty,
      eop_in => lcd_pixel_converter_in_endofpacket,
      ready_in => lcd_pixel_converter_out_ready,
      reset_n => lcd_pixel_converter_in_reset_n,
      sop_in => lcd_pixel_converter_in_startofpacket,
      valid_in => lcd_pixel_converter_in_valid
    );


  --the_lcd_pixel_fifo_in, which is an e_instance
  the_lcd_pixel_fifo_in : lcd_pixel_fifo_in_arbitrator
    port map(
      lcd_pixel_fifo_in_data => lcd_pixel_fifo_in_data,
      lcd_pixel_fifo_in_empty => lcd_pixel_fifo_in_empty,
      lcd_pixel_fifo_in_endofpacket => lcd_pixel_fifo_in_endofpacket,
      lcd_pixel_fifo_in_ready_from_sa => lcd_pixel_fifo_in_ready_from_sa,
      lcd_pixel_fifo_in_reset_n => lcd_pixel_fifo_in_reset_n,
      lcd_pixel_fifo_in_startofpacket => lcd_pixel_fifo_in_startofpacket,
      lcd_pixel_fifo_in_valid => lcd_pixel_fifo_in_valid,
      clk => internal_sdram_phy_clk_out,
      lcd_pixel_fifo_in_ready => lcd_pixel_fifo_in_ready,
      lcd_ta_sgdma_to_fifo_out_data => lcd_ta_sgdma_to_fifo_out_data,
      lcd_ta_sgdma_to_fifo_out_empty => lcd_ta_sgdma_to_fifo_out_empty,
      lcd_ta_sgdma_to_fifo_out_endofpacket => lcd_ta_sgdma_to_fifo_out_endofpacket,
      lcd_ta_sgdma_to_fifo_out_startofpacket => lcd_ta_sgdma_to_fifo_out_startofpacket,
      lcd_ta_sgdma_to_fifo_out_valid => lcd_ta_sgdma_to_fifo_out_valid,
      reset_n => sdram_phy_clk_out_reset_n
    );


  --the_lcd_pixel_fifo_out, which is an e_instance
  the_lcd_pixel_fifo_out : lcd_pixel_fifo_out_arbitrator
    port map(
      lcd_pixel_fifo_out_ready => lcd_pixel_fifo_out_ready,
      lcd_pixel_fifo_out_reset_n => lcd_pixel_fifo_out_reset_n,
      clk => clk100MHz,
      lcd_pixel_fifo_out_data => lcd_pixel_fifo_out_data,
      lcd_pixel_fifo_out_empty => lcd_pixel_fifo_out_empty,
      lcd_pixel_fifo_out_endofpacket => lcd_pixel_fifo_out_endofpacket,
      lcd_pixel_fifo_out_startofpacket => lcd_pixel_fifo_out_startofpacket,
      lcd_pixel_fifo_out_valid => lcd_pixel_fifo_out_valid,
      lcd_ta_fifo_to_dfa_in_ready_from_sa => lcd_ta_fifo_to_dfa_in_ready_from_sa,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_pixel_fifo, which is an e_ptf_instance
  the_lcd_pixel_fifo : lcd_pixel_fifo
    port map(
      avalonst_sink_ready => lcd_pixel_fifo_in_ready,
      avalonst_source_data => lcd_pixel_fifo_out_data,
      avalonst_source_empty => lcd_pixel_fifo_out_empty,
      avalonst_source_endofpacket => lcd_pixel_fifo_out_endofpacket,
      avalonst_source_startofpacket => lcd_pixel_fifo_out_startofpacket,
      avalonst_source_valid => lcd_pixel_fifo_out_valid,
      avalonst_sink_data => lcd_pixel_fifo_in_data,
      avalonst_sink_empty => lcd_pixel_fifo_in_empty,
      avalonst_sink_endofpacket => lcd_pixel_fifo_in_endofpacket,
      avalonst_sink_startofpacket => lcd_pixel_fifo_in_startofpacket,
      avalonst_sink_valid => lcd_pixel_fifo_in_valid,
      avalonst_source_ready => lcd_pixel_fifo_out_ready,
      rdclock => clk100MHz,
      rdreset_n => lcd_pixel_fifo_out_reset_n,
      wrclock => internal_sdram_phy_clk_out,
      wrreset_n => lcd_pixel_fifo_in_reset_n
    );


  --the_lcd_sgdma_csr, which is an e_instance
  the_lcd_sgdma_csr : lcd_sgdma_csr_arbitrator
    port map(
      cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr => cpu_ddr_clock_bridge_m1_granted_lcd_sgdma_csr,
      cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr => cpu_ddr_clock_bridge_m1_qualified_request_lcd_sgdma_csr,
      cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr => cpu_ddr_clock_bridge_m1_read_data_valid_lcd_sgdma_csr,
      cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr => cpu_ddr_clock_bridge_m1_requests_lcd_sgdma_csr,
      d1_lcd_sgdma_csr_end_xfer => d1_lcd_sgdma_csr_end_xfer,
      lcd_sgdma_csr_address => lcd_sgdma_csr_address,
      lcd_sgdma_csr_chipselect => lcd_sgdma_csr_chipselect,
      lcd_sgdma_csr_irq_from_sa => lcd_sgdma_csr_irq_from_sa,
      lcd_sgdma_csr_read => lcd_sgdma_csr_read,
      lcd_sgdma_csr_readdata_from_sa => lcd_sgdma_csr_readdata_from_sa,
      lcd_sgdma_csr_reset_n => lcd_sgdma_csr_reset_n,
      lcd_sgdma_csr_write => lcd_sgdma_csr_write,
      lcd_sgdma_csr_writedata => lcd_sgdma_csr_writedata,
      clk => internal_sdram_phy_clk_out,
      cpu_ddr_clock_bridge_m1_address_to_slave => cpu_ddr_clock_bridge_m1_address_to_slave,
      cpu_ddr_clock_bridge_m1_latency_counter => cpu_ddr_clock_bridge_m1_latency_counter,
      cpu_ddr_clock_bridge_m1_read => cpu_ddr_clock_bridge_m1_read,
      cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register => cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register,
      cpu_ddr_clock_bridge_m1_write => cpu_ddr_clock_bridge_m1_write,
      cpu_ddr_clock_bridge_m1_writedata => cpu_ddr_clock_bridge_m1_writedata,
      lcd_sgdma_csr_irq => lcd_sgdma_csr_irq,
      lcd_sgdma_csr_readdata => lcd_sgdma_csr_readdata,
      reset_n => sdram_phy_clk_out_reset_n
    );


  --the_lcd_sgdma_descriptor_read, which is an e_instance
  the_lcd_sgdma_descriptor_read : lcd_sgdma_descriptor_read_arbitrator
    port map(
      lcd_sgdma_descriptor_read_address_to_slave => lcd_sgdma_descriptor_read_address_to_slave,
      lcd_sgdma_descriptor_read_latency_counter => lcd_sgdma_descriptor_read_latency_counter,
      lcd_sgdma_descriptor_read_readdata => lcd_sgdma_descriptor_read_readdata,
      lcd_sgdma_descriptor_read_readdatavalid => lcd_sgdma_descriptor_read_readdatavalid,
      lcd_sgdma_descriptor_read_waitrequest => lcd_sgdma_descriptor_read_waitrequest,
      clk => internal_sdram_phy_clk_out,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      lcd_sgdma_descriptor_read_address => lcd_sgdma_descriptor_read_address,
      lcd_sgdma_descriptor_read_granted_sdram_s1 => lcd_sgdma_descriptor_read_granted_sdram_s1,
      lcd_sgdma_descriptor_read_qualified_request_sdram_s1 => lcd_sgdma_descriptor_read_qualified_request_sdram_s1,
      lcd_sgdma_descriptor_read_read => lcd_sgdma_descriptor_read_read,
      lcd_sgdma_descriptor_read_read_data_valid_sdram_s1 => lcd_sgdma_descriptor_read_read_data_valid_sdram_s1,
      lcd_sgdma_descriptor_read_read_data_valid_sdram_s1_shift_register => lcd_sgdma_descriptor_read_read_data_valid_sdram_s1_shift_register,
      lcd_sgdma_descriptor_read_requests_sdram_s1 => lcd_sgdma_descriptor_read_requests_sdram_s1,
      reset_n => sdram_phy_clk_out_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_n_from_sa => sdram_s1_waitrequest_n_from_sa
    );


  --the_lcd_sgdma_descriptor_write, which is an e_instance
  the_lcd_sgdma_descriptor_write : lcd_sgdma_descriptor_write_arbitrator
    port map(
      lcd_sgdma_descriptor_write_address_to_slave => lcd_sgdma_descriptor_write_address_to_slave,
      lcd_sgdma_descriptor_write_waitrequest => lcd_sgdma_descriptor_write_waitrequest,
      clk => internal_sdram_phy_clk_out,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      lcd_sgdma_descriptor_write_address => lcd_sgdma_descriptor_write_address,
      lcd_sgdma_descriptor_write_granted_sdram_s1 => lcd_sgdma_descriptor_write_granted_sdram_s1,
      lcd_sgdma_descriptor_write_qualified_request_sdram_s1 => lcd_sgdma_descriptor_write_qualified_request_sdram_s1,
      lcd_sgdma_descriptor_write_requests_sdram_s1 => lcd_sgdma_descriptor_write_requests_sdram_s1,
      lcd_sgdma_descriptor_write_write => lcd_sgdma_descriptor_write_write,
      lcd_sgdma_descriptor_write_writedata => lcd_sgdma_descriptor_write_writedata,
      reset_n => sdram_phy_clk_out_reset_n,
      sdram_s1_waitrequest_n_from_sa => sdram_s1_waitrequest_n_from_sa
    );


  --the_lcd_sgdma_m_read, which is an e_instance
  the_lcd_sgdma_m_read : lcd_sgdma_m_read_arbitrator
    port map(
      lcd_sgdma_m_read_address_to_slave => lcd_sgdma_m_read_address_to_slave,
      lcd_sgdma_m_read_latency_counter => lcd_sgdma_m_read_latency_counter,
      lcd_sgdma_m_read_readdata => lcd_sgdma_m_read_readdata,
      lcd_sgdma_m_read_readdatavalid => lcd_sgdma_m_read_readdatavalid,
      lcd_sgdma_m_read_waitrequest => lcd_sgdma_m_read_waitrequest,
      clk => internal_sdram_phy_clk_out,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      lcd_sgdma_m_read_address => lcd_sgdma_m_read_address,
      lcd_sgdma_m_read_granted_sdram_s1 => lcd_sgdma_m_read_granted_sdram_s1,
      lcd_sgdma_m_read_qualified_request_sdram_s1 => lcd_sgdma_m_read_qualified_request_sdram_s1,
      lcd_sgdma_m_read_read => lcd_sgdma_m_read_read,
      lcd_sgdma_m_read_read_data_valid_sdram_s1 => lcd_sgdma_m_read_read_data_valid_sdram_s1,
      lcd_sgdma_m_read_read_data_valid_sdram_s1_shift_register => lcd_sgdma_m_read_read_data_valid_sdram_s1_shift_register,
      lcd_sgdma_m_read_requests_sdram_s1 => lcd_sgdma_m_read_requests_sdram_s1,
      reset_n => sdram_phy_clk_out_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_n_from_sa => sdram_s1_waitrequest_n_from_sa
    );


  --the_lcd_sgdma_out, which is an e_instance
  the_lcd_sgdma_out : lcd_sgdma_out_arbitrator
    port map(
      lcd_sgdma_out_ready => lcd_sgdma_out_ready,
      clk => internal_sdram_phy_clk_out,
      lcd_sgdma_out_data => lcd_sgdma_out_data,
      lcd_sgdma_out_empty => lcd_sgdma_out_empty,
      lcd_sgdma_out_endofpacket => lcd_sgdma_out_endofpacket,
      lcd_sgdma_out_startofpacket => lcd_sgdma_out_startofpacket,
      lcd_sgdma_out_valid => lcd_sgdma_out_valid,
      lcd_ta_sgdma_to_fifo_in_ready_from_sa => lcd_ta_sgdma_to_fifo_in_ready_from_sa,
      reset_n => sdram_phy_clk_out_reset_n
    );


  --the_lcd_sgdma, which is an e_ptf_instance
  the_lcd_sgdma : lcd_sgdma
    port map(
      csr_irq => lcd_sgdma_csr_irq,
      csr_readdata => lcd_sgdma_csr_readdata,
      descriptor_read_address => lcd_sgdma_descriptor_read_address,
      descriptor_read_read => lcd_sgdma_descriptor_read_read,
      descriptor_write_address => lcd_sgdma_descriptor_write_address,
      descriptor_write_write => lcd_sgdma_descriptor_write_write,
      descriptor_write_writedata => lcd_sgdma_descriptor_write_writedata,
      m_read_address => lcd_sgdma_m_read_address,
      m_read_read => lcd_sgdma_m_read_read,
      out_data => lcd_sgdma_out_data,
      out_empty => lcd_sgdma_out_empty,
      out_endofpacket => lcd_sgdma_out_endofpacket,
      out_startofpacket => lcd_sgdma_out_startofpacket,
      out_valid => lcd_sgdma_out_valid,
      clk => internal_sdram_phy_clk_out,
      csr_address => lcd_sgdma_csr_address,
      csr_chipselect => lcd_sgdma_csr_chipselect,
      csr_read => lcd_sgdma_csr_read,
      csr_write => lcd_sgdma_csr_write,
      csr_writedata => lcd_sgdma_csr_writedata,
      descriptor_read_readdata => lcd_sgdma_descriptor_read_readdata,
      descriptor_read_readdatavalid => lcd_sgdma_descriptor_read_readdatavalid,
      descriptor_read_waitrequest => lcd_sgdma_descriptor_read_waitrequest,
      descriptor_write_waitrequest => lcd_sgdma_descriptor_write_waitrequest,
      m_read_readdata => lcd_sgdma_m_read_readdata,
      m_read_readdatavalid => lcd_sgdma_m_read_readdatavalid,
      m_read_waitrequest => lcd_sgdma_m_read_waitrequest,
      out_ready => lcd_sgdma_out_ready,
      system_reset_n => lcd_sgdma_csr_reset_n
    );


  --the_lcd_sync_generator_in, which is an e_instance
  the_lcd_sync_generator_in : lcd_sync_generator_in_arbitrator
    port map(
      lcd_sync_generator_in_data => lcd_sync_generator_in_data,
      lcd_sync_generator_in_empty => lcd_sync_generator_in_empty,
      lcd_sync_generator_in_endofpacket => lcd_sync_generator_in_endofpacket,
      lcd_sync_generator_in_ready_from_sa => lcd_sync_generator_in_ready_from_sa,
      lcd_sync_generator_in_reset_n => lcd_sync_generator_in_reset_n,
      lcd_sync_generator_in_startofpacket => lcd_sync_generator_in_startofpacket,
      lcd_sync_generator_in_valid => lcd_sync_generator_in_valid,
      clk => clk100MHz,
      lcd_24_to_8_bits_dfa_out_data => lcd_24_to_8_bits_dfa_out_data,
      lcd_24_to_8_bits_dfa_out_empty => lcd_24_to_8_bits_dfa_out_empty,
      lcd_24_to_8_bits_dfa_out_endofpacket => lcd_24_to_8_bits_dfa_out_endofpacket,
      lcd_24_to_8_bits_dfa_out_startofpacket => lcd_24_to_8_bits_dfa_out_startofpacket,
      lcd_24_to_8_bits_dfa_out_valid => lcd_24_to_8_bits_dfa_out_valid,
      lcd_sync_generator_in_ready => lcd_sync_generator_in_ready,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_sync_generator, which is an e_ptf_instance
  the_lcd_sync_generator : lcd_sync_generator
    port map(
      DEN => internal_DEN_from_the_lcd_sync_generator,
      HD => internal_HD_from_the_lcd_sync_generator,
      RGB_OUT => internal_RGB_OUT_from_the_lcd_sync_generator,
      VD => internal_VD_from_the_lcd_sync_generator,
      ready => lcd_sync_generator_in_ready,
      clk => clk100MHz,
      data => lcd_sync_generator_in_data,
      empty => lcd_sync_generator_in_empty,
      eop => lcd_sync_generator_in_endofpacket,
      reset_n => lcd_sync_generator_in_reset_n,
      sop => lcd_sync_generator_in_startofpacket,
      valid => lcd_sync_generator_in_valid
    );


  --the_lcd_ta_fifo_to_dfa_in, which is an e_instance
  the_lcd_ta_fifo_to_dfa_in : lcd_ta_fifo_to_dfa_in_arbitrator
    port map(
      lcd_ta_fifo_to_dfa_in_data => lcd_ta_fifo_to_dfa_in_data,
      lcd_ta_fifo_to_dfa_in_empty => lcd_ta_fifo_to_dfa_in_empty,
      lcd_ta_fifo_to_dfa_in_endofpacket => lcd_ta_fifo_to_dfa_in_endofpacket,
      lcd_ta_fifo_to_dfa_in_ready_from_sa => lcd_ta_fifo_to_dfa_in_ready_from_sa,
      lcd_ta_fifo_to_dfa_in_reset_n => lcd_ta_fifo_to_dfa_in_reset_n,
      lcd_ta_fifo_to_dfa_in_startofpacket => lcd_ta_fifo_to_dfa_in_startofpacket,
      lcd_ta_fifo_to_dfa_in_valid => lcd_ta_fifo_to_dfa_in_valid,
      clk => clk100MHz,
      lcd_pixel_fifo_out_data => lcd_pixel_fifo_out_data,
      lcd_pixel_fifo_out_empty => lcd_pixel_fifo_out_empty,
      lcd_pixel_fifo_out_endofpacket => lcd_pixel_fifo_out_endofpacket,
      lcd_pixel_fifo_out_startofpacket => lcd_pixel_fifo_out_startofpacket,
      lcd_pixel_fifo_out_valid => lcd_pixel_fifo_out_valid,
      lcd_ta_fifo_to_dfa_in_ready => lcd_ta_fifo_to_dfa_in_ready,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_ta_fifo_to_dfa_out, which is an e_instance
  the_lcd_ta_fifo_to_dfa_out : lcd_ta_fifo_to_dfa_out_arbitrator
    port map(
      lcd_ta_fifo_to_dfa_out_ready => lcd_ta_fifo_to_dfa_out_ready,
      clk => clk100MHz,
      lcd_64_to_32_bits_dfa_in_ready_from_sa => lcd_64_to_32_bits_dfa_in_ready_from_sa,
      lcd_ta_fifo_to_dfa_out_data => lcd_ta_fifo_to_dfa_out_data,
      lcd_ta_fifo_to_dfa_out_empty => lcd_ta_fifo_to_dfa_out_empty,
      lcd_ta_fifo_to_dfa_out_endofpacket => lcd_ta_fifo_to_dfa_out_endofpacket,
      lcd_ta_fifo_to_dfa_out_startofpacket => lcd_ta_fifo_to_dfa_out_startofpacket,
      lcd_ta_fifo_to_dfa_out_valid => lcd_ta_fifo_to_dfa_out_valid,
      reset_n => clk100MHz_reset_n
    );


  --the_lcd_ta_fifo_to_dfa, which is an e_ptf_instance
  the_lcd_ta_fifo_to_dfa : lcd_ta_fifo_to_dfa
    port map(
      in_ready => lcd_ta_fifo_to_dfa_in_ready,
      out_data => lcd_ta_fifo_to_dfa_out_data,
      out_empty => lcd_ta_fifo_to_dfa_out_empty,
      out_endofpacket => lcd_ta_fifo_to_dfa_out_endofpacket,
      out_startofpacket => lcd_ta_fifo_to_dfa_out_startofpacket,
      out_valid => lcd_ta_fifo_to_dfa_out_valid,
      clk => clk100MHz,
      in_data => lcd_ta_fifo_to_dfa_in_data,
      in_empty => lcd_ta_fifo_to_dfa_in_empty,
      in_endofpacket => lcd_ta_fifo_to_dfa_in_endofpacket,
      in_startofpacket => lcd_ta_fifo_to_dfa_in_startofpacket,
      in_valid => lcd_ta_fifo_to_dfa_in_valid,
      out_ready => lcd_ta_fifo_to_dfa_out_ready,
      reset_n => lcd_ta_fifo_to_dfa_in_reset_n
    );


  --the_lcd_ta_sgdma_to_fifo_in, which is an e_instance
  the_lcd_ta_sgdma_to_fifo_in : lcd_ta_sgdma_to_fifo_in_arbitrator
    port map(
      lcd_ta_sgdma_to_fifo_in_data => lcd_ta_sgdma_to_fifo_in_data,
      lcd_ta_sgdma_to_fifo_in_empty => lcd_ta_sgdma_to_fifo_in_empty,
      lcd_ta_sgdma_to_fifo_in_endofpacket => lcd_ta_sgdma_to_fifo_in_endofpacket,
      lcd_ta_sgdma_to_fifo_in_ready_from_sa => lcd_ta_sgdma_to_fifo_in_ready_from_sa,
      lcd_ta_sgdma_to_fifo_in_reset_n => lcd_ta_sgdma_to_fifo_in_reset_n,
      lcd_ta_sgdma_to_fifo_in_startofpacket => lcd_ta_sgdma_to_fifo_in_startofpacket,
      lcd_ta_sgdma_to_fifo_in_valid => lcd_ta_sgdma_to_fifo_in_valid,
      clk => internal_sdram_phy_clk_out,
      lcd_sgdma_out_data => lcd_sgdma_out_data,
      lcd_sgdma_out_empty => lcd_sgdma_out_empty,
      lcd_sgdma_out_endofpacket => lcd_sgdma_out_endofpacket,
      lcd_sgdma_out_startofpacket => lcd_sgdma_out_startofpacket,
      lcd_sgdma_out_valid => lcd_sgdma_out_valid,
      lcd_ta_sgdma_to_fifo_in_ready => lcd_ta_sgdma_to_fifo_in_ready,
      reset_n => sdram_phy_clk_out_reset_n
    );


  --the_lcd_ta_sgdma_to_fifo_out, which is an e_instance
  the_lcd_ta_sgdma_to_fifo_out : lcd_ta_sgdma_to_fifo_out_arbitrator
    port map(
      lcd_ta_sgdma_to_fifo_out_ready => lcd_ta_sgdma_to_fifo_out_ready,
      clk => internal_sdram_phy_clk_out,
      lcd_pixel_fifo_in_ready_from_sa => lcd_pixel_fifo_in_ready_from_sa,
      lcd_ta_sgdma_to_fifo_out_data => lcd_ta_sgdma_to_fifo_out_data,
      lcd_ta_sgdma_to_fifo_out_empty => lcd_ta_sgdma_to_fifo_out_empty,
      lcd_ta_sgdma_to_fifo_out_endofpacket => lcd_ta_sgdma_to_fifo_out_endofpacket,
      lcd_ta_sgdma_to_fifo_out_startofpacket => lcd_ta_sgdma_to_fifo_out_startofpacket,
      lcd_ta_sgdma_to_fifo_out_valid => lcd_ta_sgdma_to_fifo_out_valid,
      reset_n => sdram_phy_clk_out_reset_n
    );


  --the_lcd_ta_sgdma_to_fifo, which is an e_ptf_instance
  the_lcd_ta_sgdma_to_fifo : lcd_ta_sgdma_to_fifo
    port map(
      in_ready => lcd_ta_sgdma_to_fifo_in_ready,
      out_data => lcd_ta_sgdma_to_fifo_out_data,
      out_empty => lcd_ta_sgdma_to_fifo_out_empty,
      out_endofpacket => lcd_ta_sgdma_to_fifo_out_endofpacket,
      out_startofpacket => lcd_ta_sgdma_to_fifo_out_startofpacket,
      out_valid => lcd_ta_sgdma_to_fifo_out_valid,
      clk => internal_sdram_phy_clk_out,
      in_data => lcd_ta_sgdma_to_fifo_in_data,
      in_empty => lcd_ta_sgdma_to_fifo_in_empty,
      in_endofpacket => lcd_ta_sgdma_to_fifo_in_endofpacket,
      in_startofpacket => lcd_ta_sgdma_to_fifo_in_startofpacket,
      in_valid => lcd_ta_sgdma_to_fifo_in_valid,
      out_ready => lcd_ta_sgdma_to_fifo_out_ready,
      reset_n => lcd_ta_sgdma_to_fifo_in_reset_n
    );


  --the_performance_counter_control_slave, which is an e_instance
  the_performance_counter_control_slave : performance_counter_control_slave_arbitrator
    port map(
      cpuNios_data_master_granted_performance_counter_control_slave => cpuNios_data_master_granted_performance_counter_control_slave,
      cpuNios_data_master_qualified_request_performance_counter_control_slave => cpuNios_data_master_qualified_request_performance_counter_control_slave,
      cpuNios_data_master_read_data_valid_performance_counter_control_slave => cpuNios_data_master_read_data_valid_performance_counter_control_slave,
      cpuNios_data_master_requests_performance_counter_control_slave => cpuNios_data_master_requests_performance_counter_control_slave,
      d1_performance_counter_control_slave_end_xfer => d1_performance_counter_control_slave_end_xfer,
      performance_counter_control_slave_address => performance_counter_control_slave_address,
      performance_counter_control_slave_begintransfer => performance_counter_control_slave_begintransfer,
      performance_counter_control_slave_readdata_from_sa => performance_counter_control_slave_readdata_from_sa,
      performance_counter_control_slave_reset_n => performance_counter_control_slave_reset_n,
      performance_counter_control_slave_write => performance_counter_control_slave_write,
      performance_counter_control_slave_writedata => performance_counter_control_slave_writedata,
      registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave => registered_cpuNios_data_master_read_data_valid_performance_counter_control_slave,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      performance_counter_control_slave_readdata => performance_counter_control_slave_readdata,
      reset_n => clk100MHz_reset_n
    );


  --the_performance_counter, which is an e_ptf_instance
  the_performance_counter : performance_counter
    port map(
      readdata => performance_counter_control_slave_readdata,
      address => performance_counter_control_slave_address,
      begintransfer => performance_counter_control_slave_begintransfer,
      clk => clk100MHz,
      reset_n => performance_counter_control_slave_reset_n,
      write => performance_counter_control_slave_write,
      writedata => performance_counter_control_slave_writedata
    );


  --the_sdram_s1, which is an e_instance
  the_sdram_s1 : sdram_s1_arbitrator
    port map(
      cpu_ddr_clock_bridge_m1_granted_sdram_s1 => cpu_ddr_clock_bridge_m1_granted_sdram_s1,
      cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1 => cpu_ddr_clock_bridge_m1_qualified_request_sdram_s1,
      cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1 => cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1,
      cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register => cpu_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register,
      cpu_ddr_clock_bridge_m1_requests_sdram_s1 => cpu_ddr_clock_bridge_m1_requests_sdram_s1,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      lcd_sgdma_descriptor_read_granted_sdram_s1 => lcd_sgdma_descriptor_read_granted_sdram_s1,
      lcd_sgdma_descriptor_read_qualified_request_sdram_s1 => lcd_sgdma_descriptor_read_qualified_request_sdram_s1,
      lcd_sgdma_descriptor_read_read_data_valid_sdram_s1 => lcd_sgdma_descriptor_read_read_data_valid_sdram_s1,
      lcd_sgdma_descriptor_read_read_data_valid_sdram_s1_shift_register => lcd_sgdma_descriptor_read_read_data_valid_sdram_s1_shift_register,
      lcd_sgdma_descriptor_read_requests_sdram_s1 => lcd_sgdma_descriptor_read_requests_sdram_s1,
      lcd_sgdma_descriptor_write_granted_sdram_s1 => lcd_sgdma_descriptor_write_granted_sdram_s1,
      lcd_sgdma_descriptor_write_qualified_request_sdram_s1 => lcd_sgdma_descriptor_write_qualified_request_sdram_s1,
      lcd_sgdma_descriptor_write_requests_sdram_s1 => lcd_sgdma_descriptor_write_requests_sdram_s1,
      lcd_sgdma_m_read_granted_sdram_s1 => lcd_sgdma_m_read_granted_sdram_s1,
      lcd_sgdma_m_read_qualified_request_sdram_s1 => lcd_sgdma_m_read_qualified_request_sdram_s1,
      lcd_sgdma_m_read_read_data_valid_sdram_s1 => lcd_sgdma_m_read_read_data_valid_sdram_s1,
      lcd_sgdma_m_read_read_data_valid_sdram_s1_shift_register => lcd_sgdma_m_read_read_data_valid_sdram_s1_shift_register,
      lcd_sgdma_m_read_requests_sdram_s1 => lcd_sgdma_m_read_requests_sdram_s1,
      sdram_s1_address => sdram_s1_address,
      sdram_s1_beginbursttransfer => sdram_s1_beginbursttransfer,
      sdram_s1_burstcount => sdram_s1_burstcount,
      sdram_s1_byteenable => sdram_s1_byteenable,
      sdram_s1_read => sdram_s1_read,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_resetrequest_n_from_sa => sdram_s1_resetrequest_n_from_sa,
      sdram_s1_waitrequest_n_from_sa => sdram_s1_waitrequest_n_from_sa,
      sdram_s1_write => sdram_s1_write,
      sdram_s1_writedata => sdram_s1_writedata,
      tse_ddr_clock_bridge_m1_granted_sdram_s1 => tse_ddr_clock_bridge_m1_granted_sdram_s1,
      tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 => tse_ddr_clock_bridge_m1_qualified_request_sdram_s1,
      tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1 => tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1,
      tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register => tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register,
      tse_ddr_clock_bridge_m1_requests_sdram_s1 => tse_ddr_clock_bridge_m1_requests_sdram_s1,
      clk => internal_sdram_phy_clk_out,
      cpu_ddr_clock_bridge_m1_address_to_slave => cpu_ddr_clock_bridge_m1_address_to_slave,
      cpu_ddr_clock_bridge_m1_byteenable => cpu_ddr_clock_bridge_m1_byteenable,
      cpu_ddr_clock_bridge_m1_latency_counter => cpu_ddr_clock_bridge_m1_latency_counter,
      cpu_ddr_clock_bridge_m1_read => cpu_ddr_clock_bridge_m1_read,
      cpu_ddr_clock_bridge_m1_write => cpu_ddr_clock_bridge_m1_write,
      cpu_ddr_clock_bridge_m1_writedata => cpu_ddr_clock_bridge_m1_writedata,
      lcd_sgdma_descriptor_read_address_to_slave => lcd_sgdma_descriptor_read_address_to_slave,
      lcd_sgdma_descriptor_read_latency_counter => lcd_sgdma_descriptor_read_latency_counter,
      lcd_sgdma_descriptor_read_read => lcd_sgdma_descriptor_read_read,
      lcd_sgdma_descriptor_write_address_to_slave => lcd_sgdma_descriptor_write_address_to_slave,
      lcd_sgdma_descriptor_write_write => lcd_sgdma_descriptor_write_write,
      lcd_sgdma_descriptor_write_writedata => lcd_sgdma_descriptor_write_writedata,
      lcd_sgdma_m_read_address_to_slave => lcd_sgdma_m_read_address_to_slave,
      lcd_sgdma_m_read_latency_counter => lcd_sgdma_m_read_latency_counter,
      lcd_sgdma_m_read_read => lcd_sgdma_m_read_read,
      reset_n => sdram_phy_clk_out_reset_n,
      sdram_s1_readdata => sdram_s1_readdata,
      sdram_s1_readdatavalid => sdram_s1_readdatavalid,
      sdram_s1_resetrequest_n => sdram_s1_resetrequest_n,
      sdram_s1_waitrequest_n => sdram_s1_waitrequest_n,
      tse_ddr_clock_bridge_m1_address_to_slave => tse_ddr_clock_bridge_m1_address_to_slave,
      tse_ddr_clock_bridge_m1_byteenable => tse_ddr_clock_bridge_m1_byteenable,
      tse_ddr_clock_bridge_m1_latency_counter => tse_ddr_clock_bridge_m1_latency_counter,
      tse_ddr_clock_bridge_m1_read => tse_ddr_clock_bridge_m1_read,
      tse_ddr_clock_bridge_m1_write => tse_ddr_clock_bridge_m1_write,
      tse_ddr_clock_bridge_m1_writedata => tse_ddr_clock_bridge_m1_writedata
    );


  --sdram_aux_full_rate_clk_out out_clk assignment, which is an e_assign
  sdram_aux_full_rate_clk_out <= out_clk_sdram_aux_full_rate_clk;
  --sdram_aux_half_rate_clk_out out_clk assignment, which is an e_assign
  sdram_aux_half_rate_clk_out <= out_clk_sdram_aux_half_rate_clk;
  --sdram_phy_clk_out out_clk assignment, which is an e_assign
  internal_sdram_phy_clk_out <= out_clk_sdram_phy_clk;
  --reset is asserted asynchronously and deasserted synchronously
  processador_reset_clk50Mhz_domain_synch : processador_reset_clk50Mhz_domain_synch_module
    port map(
      data_out => clk50Mhz_reset_n,
      clk => clk50Mhz,
      data_in => module_input30,
      reset_n => reset_n_sources
    );

  module_input30 <= std_logic'('1');

  --reset sources mux, which is an e_mux
  reset_n_sources <= Vector_To_Std_Logic(NOT (((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT reset_n))) OR std_logic_vector'("00000000000000000000000000000000")) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpuNios_jtag_debug_module_resetrequest_from_sa)))) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_resetrequest_n_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_s1_resetrequest_n_from_sa))))));
  --the_sdram, which is an e_ptf_instance
  the_sdram : sdram
    port map(
      aux_full_rate_clk => out_clk_sdram_aux_full_rate_clk,
      aux_half_rate_clk => out_clk_sdram_aux_half_rate_clk,
      local_init_done => internal_local_init_done_from_the_sdram,
      local_rdata => sdram_s1_readdata,
      local_rdata_valid => sdram_s1_readdatavalid,
      local_ready => sdram_s1_waitrequest_n,
      local_refresh_ack => internal_local_refresh_ack_from_the_sdram,
      local_wdata_req => internal_local_wdata_req_from_the_sdram,
      mem_addr => internal_mem_addr_from_the_sdram,
      mem_ba => internal_mem_ba_from_the_sdram,
      mem_cas_n => internal_mem_cas_n_from_the_sdram,
      mem_cke(0) => internal_mem_cke_from_the_sdram,
      mem_clk(0) => mem_clk_to_and_from_the_sdram,
      mem_clk_n(0) => mem_clk_n_to_and_from_the_sdram,
      mem_cs_n(0) => internal_mem_cs_n_from_the_sdram,
      mem_dm => internal_mem_dm_from_the_sdram,
      mem_dq => mem_dq_to_and_from_the_sdram,
      mem_dqs => mem_dqs_to_and_from_the_sdram,
      mem_ras_n => internal_mem_ras_n_from_the_sdram,
      mem_we_n => internal_mem_we_n_from_the_sdram,
      phy_clk => out_clk_sdram_phy_clk,
      reset_phy_clk_n => internal_reset_phy_clk_n_from_the_sdram,
      reset_request_n => sdram_s1_resetrequest_n,
      global_reset_n => global_reset_n_to_the_sdram,
      local_address => sdram_s1_address,
      local_be => sdram_s1_byteenable,
      local_burstbegin => sdram_s1_beginbursttransfer,
      local_read_req => sdram_s1_read,
      local_size => sdram_s1_burstcount,
      local_wdata => sdram_s1_writedata,
      local_write_req => sdram_s1_write,
      pll_ref_clk => clk50Mhz,
      soft_reset_n => clk50Mhz_reset_n
    );


  --the_sgdma_rx_csr, which is an e_instance
  the_sgdma_rx_csr : sgdma_rx_csr_arbitrator
    port map(
      cpuNios_data_master_granted_sgdma_rx_csr => cpuNios_data_master_granted_sgdma_rx_csr,
      cpuNios_data_master_qualified_request_sgdma_rx_csr => cpuNios_data_master_qualified_request_sgdma_rx_csr,
      cpuNios_data_master_read_data_valid_sgdma_rx_csr => cpuNios_data_master_read_data_valid_sgdma_rx_csr,
      cpuNios_data_master_requests_sgdma_rx_csr => cpuNios_data_master_requests_sgdma_rx_csr,
      d1_sgdma_rx_csr_end_xfer => d1_sgdma_rx_csr_end_xfer,
      sgdma_rx_csr_address => sgdma_rx_csr_address,
      sgdma_rx_csr_chipselect => sgdma_rx_csr_chipselect,
      sgdma_rx_csr_irq_from_sa => sgdma_rx_csr_irq_from_sa,
      sgdma_rx_csr_read => sgdma_rx_csr_read,
      sgdma_rx_csr_readdata_from_sa => sgdma_rx_csr_readdata_from_sa,
      sgdma_rx_csr_reset_n => sgdma_rx_csr_reset_n,
      sgdma_rx_csr_write => sgdma_rx_csr_write,
      sgdma_rx_csr_writedata => sgdma_rx_csr_writedata,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      reset_n => clk100MHz_reset_n,
      sgdma_rx_csr_irq => sgdma_rx_csr_irq,
      sgdma_rx_csr_readdata => sgdma_rx_csr_readdata
    );


  --the_sgdma_rx_in, which is an e_instance
  the_sgdma_rx_in : sgdma_rx_in_arbitrator
    port map(
      sgdma_rx_in_data => sgdma_rx_in_data,
      sgdma_rx_in_empty => sgdma_rx_in_empty,
      sgdma_rx_in_endofpacket => sgdma_rx_in_endofpacket,
      sgdma_rx_in_error => sgdma_rx_in_error,
      sgdma_rx_in_ready_from_sa => sgdma_rx_in_ready_from_sa,
      sgdma_rx_in_startofpacket => sgdma_rx_in_startofpacket,
      sgdma_rx_in_valid => sgdma_rx_in_valid,
      clk => clk100MHz,
      reset_n => clk100MHz_reset_n,
      sgdma_rx_in_ready => sgdma_rx_in_ready,
      tse_mac_receive_data => tse_mac_receive_data,
      tse_mac_receive_empty => tse_mac_receive_empty,
      tse_mac_receive_endofpacket => tse_mac_receive_endofpacket,
      tse_mac_receive_error => tse_mac_receive_error,
      tse_mac_receive_startofpacket => tse_mac_receive_startofpacket,
      tse_mac_receive_valid => tse_mac_receive_valid
    );


  --the_sgdma_rx_descriptor_read, which is an e_instance
  the_sgdma_rx_descriptor_read : sgdma_rx_descriptor_read_arbitrator
    port map(
      sgdma_rx_descriptor_read_address_to_slave => sgdma_rx_descriptor_read_address_to_slave,
      sgdma_rx_descriptor_read_latency_counter => sgdma_rx_descriptor_read_latency_counter,
      sgdma_rx_descriptor_read_readdata => sgdma_rx_descriptor_read_readdata,
      sgdma_rx_descriptor_read_readdatavalid => sgdma_rx_descriptor_read_readdatavalid,
      sgdma_rx_descriptor_read_waitrequest => sgdma_rx_descriptor_read_waitrequest,
      clk => clk100MHz,
      d1_descriptor_offset_bridge_s1_end_xfer => d1_descriptor_offset_bridge_s1_end_xfer,
      descriptor_offset_bridge_s1_readdata_from_sa => descriptor_offset_bridge_s1_readdata_from_sa,
      descriptor_offset_bridge_s1_waitrequest_from_sa => descriptor_offset_bridge_s1_waitrequest_from_sa,
      reset_n => clk100MHz_reset_n,
      sgdma_rx_descriptor_read_address => sgdma_rx_descriptor_read_address,
      sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_read_granted_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_read_qualified_request_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_read_read => sgdma_rx_descriptor_read_read,
      sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register => sgdma_rx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register,
      sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_read_requests_descriptor_offset_bridge_s1
    );


  --the_sgdma_rx_descriptor_write, which is an e_instance
  the_sgdma_rx_descriptor_write : sgdma_rx_descriptor_write_arbitrator
    port map(
      sgdma_rx_descriptor_write_address_to_slave => sgdma_rx_descriptor_write_address_to_slave,
      sgdma_rx_descriptor_write_waitrequest => sgdma_rx_descriptor_write_waitrequest,
      clk => clk100MHz,
      d1_descriptor_offset_bridge_s1_end_xfer => d1_descriptor_offset_bridge_s1_end_xfer,
      descriptor_offset_bridge_s1_waitrequest_from_sa => descriptor_offset_bridge_s1_waitrequest_from_sa,
      reset_n => clk100MHz_reset_n,
      sgdma_rx_descriptor_write_address => sgdma_rx_descriptor_write_address,
      sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_write_granted_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_write_qualified_request_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1 => sgdma_rx_descriptor_write_requests_descriptor_offset_bridge_s1,
      sgdma_rx_descriptor_write_write => sgdma_rx_descriptor_write_write,
      sgdma_rx_descriptor_write_writedata => sgdma_rx_descriptor_write_writedata
    );


  --the_sgdma_rx_m_write, which is an e_instance
  the_sgdma_rx_m_write : sgdma_rx_m_write_arbitrator
    port map(
      sgdma_rx_m_write_address_to_slave => sgdma_rx_m_write_address_to_slave,
      sgdma_rx_m_write_waitrequest => sgdma_rx_m_write_waitrequest,
      clk => clk100MHz,
      d1_tse_ddr_clock_bridge_s1_end_xfer => d1_tse_ddr_clock_bridge_s1_end_xfer,
      reset_n => clk100MHz_reset_n,
      sgdma_rx_m_write_address => sgdma_rx_m_write_address,
      sgdma_rx_m_write_byteenable => sgdma_rx_m_write_byteenable,
      sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 => sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1,
      sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 => sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1,
      sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 => sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1,
      sgdma_rx_m_write_write => sgdma_rx_m_write_write,
      sgdma_rx_m_write_writedata => sgdma_rx_m_write_writedata,
      tse_ddr_clock_bridge_s1_waitrequest_from_sa => tse_ddr_clock_bridge_s1_waitrequest_from_sa
    );


  --the_sgdma_rx, which is an e_ptf_instance
  the_sgdma_rx : sgdma_rx
    port map(
      csr_irq => sgdma_rx_csr_irq,
      csr_readdata => sgdma_rx_csr_readdata,
      descriptor_read_address => sgdma_rx_descriptor_read_address,
      descriptor_read_read => sgdma_rx_descriptor_read_read,
      descriptor_write_address => sgdma_rx_descriptor_write_address,
      descriptor_write_write => sgdma_rx_descriptor_write_write,
      descriptor_write_writedata => sgdma_rx_descriptor_write_writedata,
      in_ready => sgdma_rx_in_ready,
      m_write_address => sgdma_rx_m_write_address,
      m_write_byteenable => sgdma_rx_m_write_byteenable,
      m_write_write => sgdma_rx_m_write_write,
      m_write_writedata => sgdma_rx_m_write_writedata,
      clk => clk100MHz,
      csr_address => sgdma_rx_csr_address,
      csr_chipselect => sgdma_rx_csr_chipselect,
      csr_read => sgdma_rx_csr_read,
      csr_write => sgdma_rx_csr_write,
      csr_writedata => sgdma_rx_csr_writedata,
      descriptor_read_readdata => sgdma_rx_descriptor_read_readdata,
      descriptor_read_readdatavalid => sgdma_rx_descriptor_read_readdatavalid,
      descriptor_read_waitrequest => sgdma_rx_descriptor_read_waitrequest,
      descriptor_write_waitrequest => sgdma_rx_descriptor_write_waitrequest,
      in_data => sgdma_rx_in_data,
      in_empty => sgdma_rx_in_empty,
      in_endofpacket => sgdma_rx_in_endofpacket,
      in_error => sgdma_rx_in_error,
      in_startofpacket => sgdma_rx_in_startofpacket,
      in_valid => sgdma_rx_in_valid,
      m_write_waitrequest => sgdma_rx_m_write_waitrequest,
      system_reset_n => sgdma_rx_csr_reset_n
    );


  --the_sgdma_tx_csr, which is an e_instance
  the_sgdma_tx_csr : sgdma_tx_csr_arbitrator
    port map(
      cpuNios_data_master_granted_sgdma_tx_csr => cpuNios_data_master_granted_sgdma_tx_csr,
      cpuNios_data_master_qualified_request_sgdma_tx_csr => cpuNios_data_master_qualified_request_sgdma_tx_csr,
      cpuNios_data_master_read_data_valid_sgdma_tx_csr => cpuNios_data_master_read_data_valid_sgdma_tx_csr,
      cpuNios_data_master_requests_sgdma_tx_csr => cpuNios_data_master_requests_sgdma_tx_csr,
      d1_sgdma_tx_csr_end_xfer => d1_sgdma_tx_csr_end_xfer,
      sgdma_tx_csr_address => sgdma_tx_csr_address,
      sgdma_tx_csr_chipselect => sgdma_tx_csr_chipselect,
      sgdma_tx_csr_irq_from_sa => sgdma_tx_csr_irq_from_sa,
      sgdma_tx_csr_read => sgdma_tx_csr_read,
      sgdma_tx_csr_readdata_from_sa => sgdma_tx_csr_readdata_from_sa,
      sgdma_tx_csr_reset_n => sgdma_tx_csr_reset_n,
      sgdma_tx_csr_write => sgdma_tx_csr_write,
      sgdma_tx_csr_writedata => sgdma_tx_csr_writedata,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      reset_n => clk100MHz_reset_n,
      sgdma_tx_csr_irq => sgdma_tx_csr_irq,
      sgdma_tx_csr_readdata => sgdma_tx_csr_readdata
    );


  --the_sgdma_tx_descriptor_read, which is an e_instance
  the_sgdma_tx_descriptor_read : sgdma_tx_descriptor_read_arbitrator
    port map(
      sgdma_tx_descriptor_read_address_to_slave => sgdma_tx_descriptor_read_address_to_slave,
      sgdma_tx_descriptor_read_latency_counter => sgdma_tx_descriptor_read_latency_counter,
      sgdma_tx_descriptor_read_readdata => sgdma_tx_descriptor_read_readdata,
      sgdma_tx_descriptor_read_readdatavalid => sgdma_tx_descriptor_read_readdatavalid,
      sgdma_tx_descriptor_read_waitrequest => sgdma_tx_descriptor_read_waitrequest,
      clk => clk100MHz,
      d1_descriptor_offset_bridge_s1_end_xfer => d1_descriptor_offset_bridge_s1_end_xfer,
      descriptor_offset_bridge_s1_readdata_from_sa => descriptor_offset_bridge_s1_readdata_from_sa,
      descriptor_offset_bridge_s1_waitrequest_from_sa => descriptor_offset_bridge_s1_waitrequest_from_sa,
      reset_n => clk100MHz_reset_n,
      sgdma_tx_descriptor_read_address => sgdma_tx_descriptor_read_address,
      sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_read_granted_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_read_qualified_request_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_read_read => sgdma_tx_descriptor_read_read,
      sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register => sgdma_tx_descriptor_read_read_data_valid_descriptor_offset_bridge_s1_shift_register,
      sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_read_requests_descriptor_offset_bridge_s1
    );


  --the_sgdma_tx_descriptor_write, which is an e_instance
  the_sgdma_tx_descriptor_write : sgdma_tx_descriptor_write_arbitrator
    port map(
      sgdma_tx_descriptor_write_address_to_slave => sgdma_tx_descriptor_write_address_to_slave,
      sgdma_tx_descriptor_write_waitrequest => sgdma_tx_descriptor_write_waitrequest,
      clk => clk100MHz,
      d1_descriptor_offset_bridge_s1_end_xfer => d1_descriptor_offset_bridge_s1_end_xfer,
      descriptor_offset_bridge_s1_waitrequest_from_sa => descriptor_offset_bridge_s1_waitrequest_from_sa,
      reset_n => clk100MHz_reset_n,
      sgdma_tx_descriptor_write_address => sgdma_tx_descriptor_write_address,
      sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_write_granted_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_write_qualified_request_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1 => sgdma_tx_descriptor_write_requests_descriptor_offset_bridge_s1,
      sgdma_tx_descriptor_write_write => sgdma_tx_descriptor_write_write,
      sgdma_tx_descriptor_write_writedata => sgdma_tx_descriptor_write_writedata
    );


  --the_sgdma_tx_m_read, which is an e_instance
  the_sgdma_tx_m_read : sgdma_tx_m_read_arbitrator
    port map(
      sgdma_tx_m_read_address_to_slave => sgdma_tx_m_read_address_to_slave,
      sgdma_tx_m_read_latency_counter => sgdma_tx_m_read_latency_counter,
      sgdma_tx_m_read_readdata => sgdma_tx_m_read_readdata,
      sgdma_tx_m_read_readdatavalid => sgdma_tx_m_read_readdatavalid,
      sgdma_tx_m_read_waitrequest => sgdma_tx_m_read_waitrequest,
      clk => clk100MHz,
      d1_tse_ddr_clock_bridge_s1_end_xfer => d1_tse_ddr_clock_bridge_s1_end_xfer,
      reset_n => clk100MHz_reset_n,
      sgdma_tx_m_read_address => sgdma_tx_m_read_address,
      sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 => sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1,
      sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 => sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1,
      sgdma_tx_m_read_read => sgdma_tx_m_read_read,
      sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1 => sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1,
      sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1_shift_register => sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1_shift_register,
      sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 => sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1,
      tse_ddr_clock_bridge_s1_readdata_from_sa => tse_ddr_clock_bridge_s1_readdata_from_sa,
      tse_ddr_clock_bridge_s1_waitrequest_from_sa => tse_ddr_clock_bridge_s1_waitrequest_from_sa
    );


  --the_sgdma_tx_out, which is an e_instance
  the_sgdma_tx_out : sgdma_tx_out_arbitrator
    port map(
      sgdma_tx_out_ready => sgdma_tx_out_ready,
      clk => clk100MHz,
      reset_n => clk100MHz_reset_n,
      sgdma_tx_out_data => sgdma_tx_out_data,
      sgdma_tx_out_empty => sgdma_tx_out_empty,
      sgdma_tx_out_endofpacket => sgdma_tx_out_endofpacket,
      sgdma_tx_out_error => sgdma_tx_out_error,
      sgdma_tx_out_startofpacket => sgdma_tx_out_startofpacket,
      sgdma_tx_out_valid => sgdma_tx_out_valid,
      tse_mac_transmit_ready_from_sa => tse_mac_transmit_ready_from_sa
    );


  --the_sgdma_tx, which is an e_ptf_instance
  the_sgdma_tx : sgdma_tx
    port map(
      csr_irq => sgdma_tx_csr_irq,
      csr_readdata => sgdma_tx_csr_readdata,
      descriptor_read_address => sgdma_tx_descriptor_read_address,
      descriptor_read_read => sgdma_tx_descriptor_read_read,
      descriptor_write_address => sgdma_tx_descriptor_write_address,
      descriptor_write_write => sgdma_tx_descriptor_write_write,
      descriptor_write_writedata => sgdma_tx_descriptor_write_writedata,
      m_read_address => sgdma_tx_m_read_address,
      m_read_read => sgdma_tx_m_read_read,
      out_data => sgdma_tx_out_data,
      out_empty => sgdma_tx_out_empty,
      out_endofpacket => sgdma_tx_out_endofpacket,
      out_error => sgdma_tx_out_error,
      out_startofpacket => sgdma_tx_out_startofpacket,
      out_valid => sgdma_tx_out_valid,
      clk => clk100MHz,
      csr_address => sgdma_tx_csr_address,
      csr_chipselect => sgdma_tx_csr_chipselect,
      csr_read => sgdma_tx_csr_read,
      csr_write => sgdma_tx_csr_write,
      csr_writedata => sgdma_tx_csr_writedata,
      descriptor_read_readdata => sgdma_tx_descriptor_read_readdata,
      descriptor_read_readdatavalid => sgdma_tx_descriptor_read_readdatavalid,
      descriptor_read_waitrequest => sgdma_tx_descriptor_read_waitrequest,
      descriptor_write_waitrequest => sgdma_tx_descriptor_write_waitrequest,
      m_read_readdata => sgdma_tx_m_read_readdata,
      m_read_readdatavalid => sgdma_tx_m_read_readdatavalid,
      m_read_waitrequest => sgdma_tx_m_read_waitrequest,
      out_ready => sgdma_tx_out_ready,
      system_reset_n => sgdma_tx_csr_reset_n
    );


  --the_sys_clk_timer_s1, which is an e_instance
  the_sys_clk_timer_s1 : sys_clk_timer_s1_arbitrator
    port map(
      cpuNios_data_master_granted_sys_clk_timer_s1 => cpuNios_data_master_granted_sys_clk_timer_s1,
      cpuNios_data_master_qualified_request_sys_clk_timer_s1 => cpuNios_data_master_qualified_request_sys_clk_timer_s1,
      cpuNios_data_master_read_data_valid_sys_clk_timer_s1 => cpuNios_data_master_read_data_valid_sys_clk_timer_s1,
      cpuNios_data_master_requests_sys_clk_timer_s1 => cpuNios_data_master_requests_sys_clk_timer_s1,
      d1_sys_clk_timer_s1_end_xfer => d1_sys_clk_timer_s1_end_xfer,
      sys_clk_timer_s1_address => sys_clk_timer_s1_address,
      sys_clk_timer_s1_chipselect => sys_clk_timer_s1_chipselect,
      sys_clk_timer_s1_irq_from_sa => sys_clk_timer_s1_irq_from_sa,
      sys_clk_timer_s1_readdata_from_sa => sys_clk_timer_s1_readdata_from_sa,
      sys_clk_timer_s1_reset_n => sys_clk_timer_s1_reset_n,
      sys_clk_timer_s1_write_n => sys_clk_timer_s1_write_n,
      sys_clk_timer_s1_writedata => sys_clk_timer_s1_writedata,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      reset_n => clk100MHz_reset_n,
      sys_clk_timer_s1_irq => sys_clk_timer_s1_irq,
      sys_clk_timer_s1_readdata => sys_clk_timer_s1_readdata
    );


  --the_sys_clk_timer, which is an e_ptf_instance
  the_sys_clk_timer : sys_clk_timer
    port map(
      irq => sys_clk_timer_s1_irq,
      readdata => sys_clk_timer_s1_readdata,
      address => sys_clk_timer_s1_address,
      chipselect => sys_clk_timer_s1_chipselect,
      clk => clk100MHz,
      reset_n => sys_clk_timer_s1_reset_n,
      write_n => sys_clk_timer_s1_write_n,
      writedata => sys_clk_timer_s1_writedata
    );


  --the_sysid_control_slave, which is an e_instance
  the_sysid_control_slave : sysid_control_slave_arbitrator
    port map(
      cpuNios_data_master_granted_sysid_control_slave => cpuNios_data_master_granted_sysid_control_slave,
      cpuNios_data_master_qualified_request_sysid_control_slave => cpuNios_data_master_qualified_request_sysid_control_slave,
      cpuNios_data_master_read_data_valid_sysid_control_slave => cpuNios_data_master_read_data_valid_sysid_control_slave,
      cpuNios_data_master_requests_sysid_control_slave => cpuNios_data_master_requests_sysid_control_slave,
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      sysid_control_slave_address => sysid_control_slave_address,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa,
      sysid_control_slave_reset_n => sysid_control_slave_reset_n,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_write => cpuNios_data_master_write,
      reset_n => clk100MHz_reset_n,
      sysid_control_slave_readdata => sysid_control_slave_readdata
    );


  --the_sysid, which is an e_ptf_instance
  the_sysid : sysid
    port map(
      readdata => sysid_control_slave_readdata,
      address => sysid_control_slave_address,
      clock => sysid_control_slave_clock,
      reset_n => sysid_control_slave_reset_n
    );


  --the_tse_ddr_clock_bridge_s1, which is an e_instance
  the_tse_ddr_clock_bridge_s1 : tse_ddr_clock_bridge_s1_arbitrator
    port map(
      d1_tse_ddr_clock_bridge_s1_end_xfer => d1_tse_ddr_clock_bridge_s1_end_xfer,
      sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1 => sgdma_rx_m_write_granted_tse_ddr_clock_bridge_s1,
      sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1 => sgdma_rx_m_write_qualified_request_tse_ddr_clock_bridge_s1,
      sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1 => sgdma_rx_m_write_requests_tse_ddr_clock_bridge_s1,
      sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1 => sgdma_tx_m_read_granted_tse_ddr_clock_bridge_s1,
      sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1 => sgdma_tx_m_read_qualified_request_tse_ddr_clock_bridge_s1,
      sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1 => sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1,
      sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1_shift_register => sgdma_tx_m_read_read_data_valid_tse_ddr_clock_bridge_s1_shift_register,
      sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1 => sgdma_tx_m_read_requests_tse_ddr_clock_bridge_s1,
      tse_ddr_clock_bridge_s1_address => tse_ddr_clock_bridge_s1_address,
      tse_ddr_clock_bridge_s1_byteenable => tse_ddr_clock_bridge_s1_byteenable,
      tse_ddr_clock_bridge_s1_endofpacket_from_sa => tse_ddr_clock_bridge_s1_endofpacket_from_sa,
      tse_ddr_clock_bridge_s1_nativeaddress => tse_ddr_clock_bridge_s1_nativeaddress,
      tse_ddr_clock_bridge_s1_read => tse_ddr_clock_bridge_s1_read,
      tse_ddr_clock_bridge_s1_readdata_from_sa => tse_ddr_clock_bridge_s1_readdata_from_sa,
      tse_ddr_clock_bridge_s1_reset_n => tse_ddr_clock_bridge_s1_reset_n,
      tse_ddr_clock_bridge_s1_waitrequest_from_sa => tse_ddr_clock_bridge_s1_waitrequest_from_sa,
      tse_ddr_clock_bridge_s1_write => tse_ddr_clock_bridge_s1_write,
      tse_ddr_clock_bridge_s1_writedata => tse_ddr_clock_bridge_s1_writedata,
      clk => clk100MHz,
      reset_n => clk100MHz_reset_n,
      sgdma_rx_m_write_address_to_slave => sgdma_rx_m_write_address_to_slave,
      sgdma_rx_m_write_byteenable => sgdma_rx_m_write_byteenable,
      sgdma_rx_m_write_write => sgdma_rx_m_write_write,
      sgdma_rx_m_write_writedata => sgdma_rx_m_write_writedata,
      sgdma_tx_m_read_address_to_slave => sgdma_tx_m_read_address_to_slave,
      sgdma_tx_m_read_latency_counter => sgdma_tx_m_read_latency_counter,
      sgdma_tx_m_read_read => sgdma_tx_m_read_read,
      tse_ddr_clock_bridge_s1_endofpacket => tse_ddr_clock_bridge_s1_endofpacket,
      tse_ddr_clock_bridge_s1_readdata => tse_ddr_clock_bridge_s1_readdata,
      tse_ddr_clock_bridge_s1_readdatavalid => tse_ddr_clock_bridge_s1_readdatavalid,
      tse_ddr_clock_bridge_s1_waitrequest => tse_ddr_clock_bridge_s1_waitrequest
    );


  --the_tse_ddr_clock_bridge_m1, which is an e_instance
  the_tse_ddr_clock_bridge_m1 : tse_ddr_clock_bridge_m1_arbitrator
    port map(
      tse_ddr_clock_bridge_m1_address_to_slave => tse_ddr_clock_bridge_m1_address_to_slave,
      tse_ddr_clock_bridge_m1_latency_counter => tse_ddr_clock_bridge_m1_latency_counter,
      tse_ddr_clock_bridge_m1_readdata => tse_ddr_clock_bridge_m1_readdata,
      tse_ddr_clock_bridge_m1_readdatavalid => tse_ddr_clock_bridge_m1_readdatavalid,
      tse_ddr_clock_bridge_m1_reset_n => tse_ddr_clock_bridge_m1_reset_n,
      tse_ddr_clock_bridge_m1_waitrequest => tse_ddr_clock_bridge_m1_waitrequest,
      clk => internal_sdram_phy_clk_out,
      d1_sdram_s1_end_xfer => d1_sdram_s1_end_xfer,
      reset_n => sdram_phy_clk_out_reset_n,
      sdram_s1_readdata_from_sa => sdram_s1_readdata_from_sa,
      sdram_s1_waitrequest_n_from_sa => sdram_s1_waitrequest_n_from_sa,
      tse_ddr_clock_bridge_m1_address => tse_ddr_clock_bridge_m1_address,
      tse_ddr_clock_bridge_m1_byteenable => tse_ddr_clock_bridge_m1_byteenable,
      tse_ddr_clock_bridge_m1_granted_sdram_s1 => tse_ddr_clock_bridge_m1_granted_sdram_s1,
      tse_ddr_clock_bridge_m1_qualified_request_sdram_s1 => tse_ddr_clock_bridge_m1_qualified_request_sdram_s1,
      tse_ddr_clock_bridge_m1_read => tse_ddr_clock_bridge_m1_read,
      tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1 => tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1,
      tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register => tse_ddr_clock_bridge_m1_read_data_valid_sdram_s1_shift_register,
      tse_ddr_clock_bridge_m1_requests_sdram_s1 => tse_ddr_clock_bridge_m1_requests_sdram_s1,
      tse_ddr_clock_bridge_m1_write => tse_ddr_clock_bridge_m1_write,
      tse_ddr_clock_bridge_m1_writedata => tse_ddr_clock_bridge_m1_writedata
    );


  --the_tse_ddr_clock_bridge, which is an e_ptf_instance
  the_tse_ddr_clock_bridge : tse_ddr_clock_bridge
    port map(
      master_address => tse_ddr_clock_bridge_m1_address,
      master_byteenable => tse_ddr_clock_bridge_m1_byteenable,
      master_nativeaddress => tse_ddr_clock_bridge_m1_nativeaddress,
      master_read => tse_ddr_clock_bridge_m1_read,
      master_write => tse_ddr_clock_bridge_m1_write,
      master_writedata => tse_ddr_clock_bridge_m1_writedata,
      slave_endofpacket => tse_ddr_clock_bridge_s1_endofpacket,
      slave_readdata => tse_ddr_clock_bridge_s1_readdata,
      slave_readdatavalid => tse_ddr_clock_bridge_s1_readdatavalid,
      slave_waitrequest => tse_ddr_clock_bridge_s1_waitrequest,
      master_clk => internal_sdram_phy_clk_out,
      master_endofpacket => tse_ddr_clock_bridge_m1_endofpacket,
      master_readdata => tse_ddr_clock_bridge_m1_readdata,
      master_readdatavalid => tse_ddr_clock_bridge_m1_readdatavalid,
      master_reset_n => tse_ddr_clock_bridge_m1_reset_n,
      master_waitrequest => tse_ddr_clock_bridge_m1_waitrequest,
      slave_address => tse_ddr_clock_bridge_s1_address,
      slave_byteenable => tse_ddr_clock_bridge_s1_byteenable,
      slave_clk => clk100MHz,
      slave_nativeaddress => tse_ddr_clock_bridge_s1_nativeaddress,
      slave_read => tse_ddr_clock_bridge_s1_read,
      slave_reset_n => tse_ddr_clock_bridge_s1_reset_n,
      slave_write => tse_ddr_clock_bridge_s1_write,
      slave_writedata => tse_ddr_clock_bridge_s1_writedata
    );


  --the_tse_mac_control_port, which is an e_instance
  the_tse_mac_control_port : tse_mac_control_port_arbitrator
    port map(
      cpuNios_data_master_granted_tse_mac_control_port => cpuNios_data_master_granted_tse_mac_control_port,
      cpuNios_data_master_qualified_request_tse_mac_control_port => cpuNios_data_master_qualified_request_tse_mac_control_port,
      cpuNios_data_master_read_data_valid_tse_mac_control_port => cpuNios_data_master_read_data_valid_tse_mac_control_port,
      cpuNios_data_master_requests_tse_mac_control_port => cpuNios_data_master_requests_tse_mac_control_port,
      d1_tse_mac_control_port_end_xfer => d1_tse_mac_control_port_end_xfer,
      tse_mac_control_port_address => tse_mac_control_port_address,
      tse_mac_control_port_read => tse_mac_control_port_read,
      tse_mac_control_port_readdata_from_sa => tse_mac_control_port_readdata_from_sa,
      tse_mac_control_port_reset => tse_mac_control_port_reset,
      tse_mac_control_port_waitrequest_from_sa => tse_mac_control_port_waitrequest_from_sa,
      tse_mac_control_port_write => tse_mac_control_port_write,
      tse_mac_control_port_writedata => tse_mac_control_port_writedata,
      clk => clk100MHz,
      cpuNios_data_master_address_to_slave => cpuNios_data_master_address_to_slave,
      cpuNios_data_master_read => cpuNios_data_master_read,
      cpuNios_data_master_waitrequest => cpuNios_data_master_waitrequest,
      cpuNios_data_master_write => cpuNios_data_master_write,
      cpuNios_data_master_writedata => cpuNios_data_master_writedata,
      reset_n => clk100MHz_reset_n,
      tse_mac_control_port_readdata => tse_mac_control_port_readdata,
      tse_mac_control_port_waitrequest => tse_mac_control_port_waitrequest
    );


  --the_tse_mac_transmit, which is an e_instance
  the_tse_mac_transmit : tse_mac_transmit_arbitrator
    port map(
      tse_mac_transmit_data => tse_mac_transmit_data,
      tse_mac_transmit_empty => tse_mac_transmit_empty,
      tse_mac_transmit_endofpacket => tse_mac_transmit_endofpacket,
      tse_mac_transmit_error => tse_mac_transmit_error,
      tse_mac_transmit_ready_from_sa => tse_mac_transmit_ready_from_sa,
      tse_mac_transmit_startofpacket => tse_mac_transmit_startofpacket,
      tse_mac_transmit_valid => tse_mac_transmit_valid,
      clk => clk100MHz,
      reset_n => clk100MHz_reset_n,
      sgdma_tx_out_data => sgdma_tx_out_data,
      sgdma_tx_out_empty => sgdma_tx_out_empty,
      sgdma_tx_out_endofpacket => sgdma_tx_out_endofpacket,
      sgdma_tx_out_error => sgdma_tx_out_error,
      sgdma_tx_out_startofpacket => sgdma_tx_out_startofpacket,
      sgdma_tx_out_valid => sgdma_tx_out_valid,
      tse_mac_transmit_ready => tse_mac_transmit_ready
    );


  --the_tse_mac_receive, which is an e_instance
  the_tse_mac_receive : tse_mac_receive_arbitrator
    port map(
      tse_mac_receive_ready => tse_mac_receive_ready,
      clk => clk100MHz,
      reset_n => clk100MHz_reset_n,
      sgdma_rx_in_ready_from_sa => sgdma_rx_in_ready_from_sa,
      tse_mac_receive_data => tse_mac_receive_data,
      tse_mac_receive_empty => tse_mac_receive_empty,
      tse_mac_receive_endofpacket => tse_mac_receive_endofpacket,
      tse_mac_receive_error => tse_mac_receive_error,
      tse_mac_receive_startofpacket => tse_mac_receive_startofpacket,
      tse_mac_receive_valid => tse_mac_receive_valid
    );


  --the_tse_mac, which is an e_ptf_instance
  the_tse_mac : tse_mac
    port map(
      ena_10 => internal_ena_10_from_the_tse_mac,
      eth_mode => internal_eth_mode_from_the_tse_mac,
      ff_rx_data => tse_mac_receive_data,
      ff_rx_dval => tse_mac_receive_valid,
      ff_rx_eop => tse_mac_receive_endofpacket,
      ff_rx_mod => tse_mac_receive_empty,
      ff_rx_sop => tse_mac_receive_startofpacket,
      ff_tx_rdy => tse_mac_transmit_ready,
      gm_tx_d => internal_gm_tx_d_from_the_tse_mac,
      gm_tx_en => internal_gm_tx_en_from_the_tse_mac,
      gm_tx_err => internal_gm_tx_err_from_the_tse_mac,
      m_tx_d => internal_m_tx_d_from_the_tse_mac,
      m_tx_en => internal_m_tx_en_from_the_tse_mac,
      m_tx_err => internal_m_tx_err_from_the_tse_mac,
      mdc => internal_mdc_from_the_tse_mac,
      mdio_oen => internal_mdio_oen_from_the_tse_mac,
      mdio_out => internal_mdio_out_from_the_tse_mac,
      readdata => tse_mac_control_port_readdata,
      rx_err => tse_mac_receive_error,
      waitrequest => tse_mac_control_port_waitrequest,
      address => tse_mac_control_port_address,
      clk => clk100MHz,
      ff_rx_clk => clk100MHz,
      ff_rx_rdy => tse_mac_receive_ready,
      ff_tx_clk => clk100MHz,
      ff_tx_data => tse_mac_transmit_data,
      ff_tx_eop => tse_mac_transmit_endofpacket,
      ff_tx_err => tse_mac_transmit_error,
      ff_tx_mod => tse_mac_transmit_empty,
      ff_tx_sop => tse_mac_transmit_startofpacket,
      ff_tx_wren => tse_mac_transmit_valid,
      gm_rx_d => gm_rx_d_to_the_tse_mac,
      gm_rx_dv => gm_rx_dv_to_the_tse_mac,
      gm_rx_err => gm_rx_err_to_the_tse_mac,
      m_rx_col => m_rx_col_to_the_tse_mac,
      m_rx_crs => m_rx_crs_to_the_tse_mac,
      m_rx_d => m_rx_d_to_the_tse_mac,
      m_rx_en => m_rx_en_to_the_tse_mac,
      m_rx_err => m_rx_err_to_the_tse_mac,
      mdio_in => mdio_in_to_the_tse_mac,
      read => tse_mac_control_port_read,
      reset => tse_mac_control_port_reset,
      rx_clk => rx_clk_to_the_tse_mac,
      set_10 => set_10_to_the_tse_mac,
      set_1000 => set_1000_to_the_tse_mac,
      tx_clk => tx_clk_to_the_tse_mac,
      write => tse_mac_control_port_write,
      writedata => tse_mac_control_port_writedata
    );


  --reset is asserted asynchronously and deasserted synchronously
  processador_reset_clk100MHz_domain_synch : processador_reset_clk100MHz_domain_synch_module
    port map(
      data_out => clk100MHz_reset_n,
      clk => clk100MHz,
      data_in => module_input43,
      reset_n => reset_n_sources
    );

  module_input43 <= std_logic'('1');

  --reset is asserted asynchronously and deasserted synchronously
  processador_reset_sdram_phy_clk_out_domain_synch : processador_reset_sdram_phy_clk_out_domain_synch_module
    port map(
      data_out => sdram_phy_clk_out_reset_n,
      clk => internal_sdram_phy_clk_out,
      data_in => module_input44,
      reset_n => reset_n_sources
    );

  module_input44 <= std_logic'('1');

  --cpu_ddr_clock_bridge_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  cpu_ddr_clock_bridge_m1_endofpacket <= std_logic'('0');
  --descriptor_offset_bridge_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  descriptor_offset_bridge_m1_endofpacket <= std_logic'('0');
  --sysid_control_slave_clock of type clock does not connect to anything so wire it to default (0)
  sysid_control_slave_clock <= std_logic'('0');
  --tse_ddr_clock_bridge_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  tse_ddr_clock_bridge_m1_endofpacket <= std_logic'('0');
  --vhdl renameroo for output signals
  DEN_from_the_lcd_sync_generator <= internal_DEN_from_the_lcd_sync_generator;
  --vhdl renameroo for output signals
  HD_from_the_lcd_sync_generator <= internal_HD_from_the_lcd_sync_generator;
  --vhdl renameroo for output signals
  RGB_OUT_from_the_lcd_sync_generator <= internal_RGB_OUT_from_the_lcd_sync_generator;
  --vhdl renameroo for output signals
  VD_from_the_lcd_sync_generator <= internal_VD_from_the_lcd_sync_generator;
  --vhdl renameroo for output signals
  counter_from_the_fft_pipeline_0 <= internal_counter_from_the_fft_pipeline_0;
  --vhdl renameroo for output signals
  ena_10_from_the_tse_mac <= internal_ena_10_from_the_tse_mac;
  --vhdl renameroo for output signals
  eth_mode_from_the_tse_mac <= internal_eth_mode_from_the_tse_mac;
  --vhdl renameroo for output signals
  gm_tx_d_from_the_tse_mac <= internal_gm_tx_d_from_the_tse_mac;
  --vhdl renameroo for output signals
  gm_tx_en_from_the_tse_mac <= internal_gm_tx_en_from_the_tse_mac;
  --vhdl renameroo for output signals
  gm_tx_err_from_the_tse_mac <= internal_gm_tx_err_from_the_tse_mac;
  --vhdl renameroo for output signals
  local_init_done_from_the_sdram <= internal_local_init_done_from_the_sdram;
  --vhdl renameroo for output signals
  local_refresh_ack_from_the_sdram <= internal_local_refresh_ack_from_the_sdram;
  --vhdl renameroo for output signals
  local_wdata_req_from_the_sdram <= internal_local_wdata_req_from_the_sdram;
  --vhdl renameroo for output signals
  m_tx_d_from_the_tse_mac <= internal_m_tx_d_from_the_tse_mac;
  --vhdl renameroo for output signals
  m_tx_en_from_the_tse_mac <= internal_m_tx_en_from_the_tse_mac;
  --vhdl renameroo for output signals
  m_tx_err_from_the_tse_mac <= internal_m_tx_err_from_the_tse_mac;
  --vhdl renameroo for output signals
  mdc_from_the_tse_mac <= internal_mdc_from_the_tse_mac;
  --vhdl renameroo for output signals
  mdio_oen_from_the_tse_mac <= internal_mdio_oen_from_the_tse_mac;
  --vhdl renameroo for output signals
  mdio_out_from_the_tse_mac <= internal_mdio_out_from_the_tse_mac;
  --vhdl renameroo for output signals
  mem_addr_from_the_sdram <= internal_mem_addr_from_the_sdram;
  --vhdl renameroo for output signals
  mem_ba_from_the_sdram <= internal_mem_ba_from_the_sdram;
  --vhdl renameroo for output signals
  mem_cas_n_from_the_sdram <= internal_mem_cas_n_from_the_sdram;
  --vhdl renameroo for output signals
  mem_cke_from_the_sdram <= internal_mem_cke_from_the_sdram;
  --vhdl renameroo for output signals
  mem_cs_n_from_the_sdram <= internal_mem_cs_n_from_the_sdram;
  --vhdl renameroo for output signals
  mem_dm_from_the_sdram <= internal_mem_dm_from_the_sdram;
  --vhdl renameroo for output signals
  mem_ras_n_from_the_sdram <= internal_mem_ras_n_from_the_sdram;
  --vhdl renameroo for output signals
  mem_we_n_from_the_sdram <= internal_mem_we_n_from_the_sdram;
  --vhdl renameroo for output signals
  out_port_from_the_lcd_i2c_en <= internal_out_port_from_the_lcd_i2c_en;
  --vhdl renameroo for output signals
  out_port_from_the_lcd_i2c_scl <= internal_out_port_from_the_lcd_i2c_scl;
  --vhdl renameroo for output signals
  reset_phy_clk_n_from_the_sdram <= internal_reset_phy_clk_n_from_the_sdram;
  --vhdl renameroo for output signals
  sdram_phy_clk_out <= internal_sdram_phy_clk_out;
  --vhdl renameroo for output signals
  tx_out_from_the_fft_pipeline_0 <= internal_tx_out_from_the_fft_pipeline_0;

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your libraries here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>

entity test_bench is 
end entity test_bench;


architecture europa of test_bench is
component processador is 
           port (
                 -- 1) global signals:
                    signal clk100MHz : IN STD_LOGIC;
                    signal clk50Mhz : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_aux_full_rate_clk_out : OUT STD_LOGIC;
                    signal sdram_aux_half_rate_clk_out : OUT STD_LOGIC;
                    signal sdram_phy_clk_out : OUT STD_LOGIC;

                 -- the_fft_pipeline_0
                    signal counter_from_the_fft_pipeline_0 : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
                    signal rx_in_to_the_fft_pipeline_0 : IN STD_LOGIC;
                    signal tx_out_from_the_fft_pipeline_0 : OUT STD_LOGIC;

                 -- the_lcd_i2c_en
                    signal out_port_from_the_lcd_i2c_en : OUT STD_LOGIC;

                 -- the_lcd_i2c_scl
                    signal out_port_from_the_lcd_i2c_scl : OUT STD_LOGIC;

                 -- the_lcd_i2c_sdat
                    signal bidir_port_to_and_from_the_lcd_i2c_sdat : INOUT STD_LOGIC;

                 -- the_lcd_sync_generator
                    signal DEN_from_the_lcd_sync_generator : OUT STD_LOGIC;
                    signal HD_from_the_lcd_sync_generator : OUT STD_LOGIC;
                    signal RGB_OUT_from_the_lcd_sync_generator : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal VD_from_the_lcd_sync_generator : OUT STD_LOGIC;

                 -- the_sdram
                    signal global_reset_n_to_the_sdram : IN STD_LOGIC;
                    signal local_init_done_from_the_sdram : OUT STD_LOGIC;
                    signal local_refresh_ack_from_the_sdram : OUT STD_LOGIC;
                    signal local_wdata_req_from_the_sdram : OUT STD_LOGIC;
                    signal mem_addr_from_the_sdram : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal mem_ba_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_cas_n_from_the_sdram : OUT STD_LOGIC;
                    signal mem_cke_from_the_sdram : OUT STD_LOGIC;
                    signal mem_clk_n_to_and_from_the_sdram : INOUT STD_LOGIC;
                    signal mem_clk_to_and_from_the_sdram : INOUT STD_LOGIC;
                    signal mem_cs_n_from_the_sdram : OUT STD_LOGIC;
                    signal mem_dm_from_the_sdram : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_dq_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal mem_dqs_to_and_from_the_sdram : INOUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal mem_ras_n_from_the_sdram : OUT STD_LOGIC;
                    signal mem_we_n_from_the_sdram : OUT STD_LOGIC;
                    signal reset_phy_clk_n_from_the_sdram : OUT STD_LOGIC;

                 -- the_tse_mac
                    signal ena_10_from_the_tse_mac : OUT STD_LOGIC;
                    signal eth_mode_from_the_tse_mac : OUT STD_LOGIC;
                    signal gm_rx_d_to_the_tse_mac : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_rx_dv_to_the_tse_mac : IN STD_LOGIC;
                    signal gm_rx_err_to_the_tse_mac : IN STD_LOGIC;
                    signal gm_tx_d_from_the_tse_mac : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_tx_en_from_the_tse_mac : OUT STD_LOGIC;
                    signal gm_tx_err_from_the_tse_mac : OUT STD_LOGIC;
                    signal m_rx_col_to_the_tse_mac : IN STD_LOGIC;
                    signal m_rx_crs_to_the_tse_mac : IN STD_LOGIC;
                    signal m_rx_d_to_the_tse_mac : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_rx_en_to_the_tse_mac : IN STD_LOGIC;
                    signal m_rx_err_to_the_tse_mac : IN STD_LOGIC;
                    signal m_tx_d_from_the_tse_mac : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_tx_en_from_the_tse_mac : OUT STD_LOGIC;
                    signal m_tx_err_from_the_tse_mac : OUT STD_LOGIC;
                    signal mdc_from_the_tse_mac : OUT STD_LOGIC;
                    signal mdio_in_to_the_tse_mac : IN STD_LOGIC;
                    signal mdio_oen_from_the_tse_mac : OUT STD_LOGIC;
                    signal mdio_out_from_the_tse_mac : OUT STD_LOGIC;
                    signal rx_clk_to_the_tse_mac : IN STD_LOGIC;
                    signal set_1000_to_the_tse_mac : IN STD_LOGIC;
                    signal set_10_to_the_tse_mac : IN STD_LOGIC;
                    signal tx_clk_to_the_tse_mac : IN STD_LOGIC
                 );
end component processador;

component tse_mac_loopback is 
           port (
                 -- inputs:
                    signal gm_tx_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_tx_en : IN STD_LOGIC;
                    signal gm_tx_err : IN STD_LOGIC;
                    signal m_tx_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_tx_en : IN STD_LOGIC;
                    signal m_tx_err : IN STD_LOGIC;

                 -- outputs:
                    signal gm_rx_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_rx_dv : OUT STD_LOGIC;
                    signal gm_rx_err : OUT STD_LOGIC;
                    signal m_rx_col : OUT STD_LOGIC;
                    signal m_rx_crs : OUT STD_LOGIC;
                    signal m_rx_d : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_rx_en : OUT STD_LOGIC;
                    signal m_rx_err : OUT STD_LOGIC;
                    signal rx_clk : OUT STD_LOGIC;
                    signal set_10 : OUT STD_LOGIC;
                    signal set_1000 : OUT STD_LOGIC;
                    signal tx_clk : OUT STD_LOGIC
                 );
end component tse_mac_loopback;

                signal DEN_from_the_lcd_sync_generator :  STD_LOGIC;
                signal HD_from_the_lcd_sync_generator :  STD_LOGIC;
                signal RGB_OUT_from_the_lcd_sync_generator :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal VD_from_the_lcd_sync_generator :  STD_LOGIC;
                signal bidir_port_to_and_from_the_lcd_i2c_sdat :  STD_LOGIC;
                signal clk :  STD_LOGIC;
                signal clk100MHz :  STD_LOGIC;
                signal clk50Mhz :  STD_LOGIC;
                signal counter_from_the_fft_pipeline_0 :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal cpu_ddr_clock_bridge_m1_endofpacket :  STD_LOGIC;
                signal cpu_ddr_clock_bridge_m1_nativeaddress :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal cpu_ddr_clock_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_debugaccess :  STD_LOGIC;
                signal descriptor_offset_bridge_m1_endofpacket :  STD_LOGIC;
                signal descriptor_offset_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal ena_10_from_the_tse_mac :  STD_LOGIC;
                signal eth_mode_from_the_tse_mac :  STD_LOGIC;
                signal global_reset_n_to_the_sdram :  STD_LOGIC;
                signal gm_rx_d_to_the_tse_mac :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gm_rx_dv_to_the_tse_mac :  STD_LOGIC;
                signal gm_rx_err_to_the_tse_mac :  STD_LOGIC;
                signal gm_tx_d_from_the_tse_mac :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gm_tx_en_from_the_tse_mac :  STD_LOGIC;
                signal gm_tx_err_from_the_tse_mac :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal local_init_done_from_the_sdram :  STD_LOGIC;
                signal local_refresh_ack_from_the_sdram :  STD_LOGIC;
                signal local_wdata_req_from_the_sdram :  STD_LOGIC;
                signal m_rx_col_to_the_tse_mac :  STD_LOGIC;
                signal m_rx_crs_to_the_tse_mac :  STD_LOGIC;
                signal m_rx_d_to_the_tse_mac :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal m_rx_en_to_the_tse_mac :  STD_LOGIC;
                signal m_rx_err_to_the_tse_mac :  STD_LOGIC;
                signal m_tx_d_from_the_tse_mac :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal m_tx_en_from_the_tse_mac :  STD_LOGIC;
                signal m_tx_err_from_the_tse_mac :  STD_LOGIC;
                signal mdc_from_the_tse_mac :  STD_LOGIC;
                signal mdio_in_to_the_tse_mac :  STD_LOGIC;
                signal mdio_oen_from_the_tse_mac :  STD_LOGIC;
                signal mdio_out_from_the_tse_mac :  STD_LOGIC;
                signal mem_addr_from_the_sdram :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal mem_ba_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal mem_cas_n_from_the_sdram :  STD_LOGIC;
                signal mem_cke_from_the_sdram :  STD_LOGIC;
                signal mem_clk_n_to_and_from_the_sdram :  STD_LOGIC;
                signal mem_clk_to_and_from_the_sdram :  STD_LOGIC;
                signal mem_cs_n_from_the_sdram :  STD_LOGIC;
                signal mem_dm_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal mem_dq_to_and_from_the_sdram :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal mem_dqs_to_and_from_the_sdram :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal mem_ras_n_from_the_sdram :  STD_LOGIC;
                signal mem_we_n_from_the_sdram :  STD_LOGIC;
                signal out_port_from_the_lcd_i2c_en :  STD_LOGIC;
                signal out_port_from_the_lcd_i2c_scl :  STD_LOGIC;
                signal reset_n :  STD_LOGIC;
                signal reset_phy_clk_n_from_the_sdram :  STD_LOGIC;
                signal rx_clk_to_the_tse_mac :  STD_LOGIC;
                signal rx_in_to_the_fft_pipeline_0 :  STD_LOGIC;
                signal sdram_aux_full_rate_clk_out :  STD_LOGIC;
                signal sdram_aux_half_rate_clk_out :  STD_LOGIC;
                signal sdram_phy_clk_out :  STD_LOGIC;
                signal set_1000_to_the_tse_mac :  STD_LOGIC;
                signal set_10_to_the_tse_mac :  STD_LOGIC;
                signal sysid_control_slave_clock :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_endofpacket :  STD_LOGIC;
                signal tse_ddr_clock_bridge_m1_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal tse_ddr_clock_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal tx_clk_to_the_tse_mac :  STD_LOGIC;
                signal tx_out_from_the_fft_pipeline_0 :  STD_LOGIC;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your component and signal declaration here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


begin

  --Set us up the Dut
  DUT : processador
    port map(
      DEN_from_the_lcd_sync_generator => DEN_from_the_lcd_sync_generator,
      HD_from_the_lcd_sync_generator => HD_from_the_lcd_sync_generator,
      RGB_OUT_from_the_lcd_sync_generator => RGB_OUT_from_the_lcd_sync_generator,
      VD_from_the_lcd_sync_generator => VD_from_the_lcd_sync_generator,
      bidir_port_to_and_from_the_lcd_i2c_sdat => bidir_port_to_and_from_the_lcd_i2c_sdat,
      counter_from_the_fft_pipeline_0 => counter_from_the_fft_pipeline_0,
      ena_10_from_the_tse_mac => ena_10_from_the_tse_mac,
      eth_mode_from_the_tse_mac => eth_mode_from_the_tse_mac,
      gm_tx_d_from_the_tse_mac => gm_tx_d_from_the_tse_mac,
      gm_tx_en_from_the_tse_mac => gm_tx_en_from_the_tse_mac,
      gm_tx_err_from_the_tse_mac => gm_tx_err_from_the_tse_mac,
      local_init_done_from_the_sdram => local_init_done_from_the_sdram,
      local_refresh_ack_from_the_sdram => local_refresh_ack_from_the_sdram,
      local_wdata_req_from_the_sdram => local_wdata_req_from_the_sdram,
      m_tx_d_from_the_tse_mac => m_tx_d_from_the_tse_mac,
      m_tx_en_from_the_tse_mac => m_tx_en_from_the_tse_mac,
      m_tx_err_from_the_tse_mac => m_tx_err_from_the_tse_mac,
      mdc_from_the_tse_mac => mdc_from_the_tse_mac,
      mdio_oen_from_the_tse_mac => mdio_oen_from_the_tse_mac,
      mdio_out_from_the_tse_mac => mdio_out_from_the_tse_mac,
      mem_addr_from_the_sdram => mem_addr_from_the_sdram,
      mem_ba_from_the_sdram => mem_ba_from_the_sdram,
      mem_cas_n_from_the_sdram => mem_cas_n_from_the_sdram,
      mem_cke_from_the_sdram => mem_cke_from_the_sdram,
      mem_clk_n_to_and_from_the_sdram => mem_clk_n_to_and_from_the_sdram,
      mem_clk_to_and_from_the_sdram => mem_clk_to_and_from_the_sdram,
      mem_cs_n_from_the_sdram => mem_cs_n_from_the_sdram,
      mem_dm_from_the_sdram => mem_dm_from_the_sdram,
      mem_dq_to_and_from_the_sdram => mem_dq_to_and_from_the_sdram,
      mem_dqs_to_and_from_the_sdram => mem_dqs_to_and_from_the_sdram,
      mem_ras_n_from_the_sdram => mem_ras_n_from_the_sdram,
      mem_we_n_from_the_sdram => mem_we_n_from_the_sdram,
      out_port_from_the_lcd_i2c_en => out_port_from_the_lcd_i2c_en,
      out_port_from_the_lcd_i2c_scl => out_port_from_the_lcd_i2c_scl,
      reset_phy_clk_n_from_the_sdram => reset_phy_clk_n_from_the_sdram,
      sdram_aux_full_rate_clk_out => sdram_aux_full_rate_clk_out,
      sdram_aux_half_rate_clk_out => sdram_aux_half_rate_clk_out,
      sdram_phy_clk_out => sdram_phy_clk_out,
      tx_out_from_the_fft_pipeline_0 => tx_out_from_the_fft_pipeline_0,
      clk100MHz => clk100MHz,
      clk50Mhz => clk50Mhz,
      global_reset_n_to_the_sdram => global_reset_n_to_the_sdram,
      gm_rx_d_to_the_tse_mac => gm_rx_d_to_the_tse_mac,
      gm_rx_dv_to_the_tse_mac => gm_rx_dv_to_the_tse_mac,
      gm_rx_err_to_the_tse_mac => gm_rx_err_to_the_tse_mac,
      m_rx_col_to_the_tse_mac => m_rx_col_to_the_tse_mac,
      m_rx_crs_to_the_tse_mac => m_rx_crs_to_the_tse_mac,
      m_rx_d_to_the_tse_mac => m_rx_d_to_the_tse_mac,
      m_rx_en_to_the_tse_mac => m_rx_en_to_the_tse_mac,
      m_rx_err_to_the_tse_mac => m_rx_err_to_the_tse_mac,
      mdio_in_to_the_tse_mac => mdio_in_to_the_tse_mac,
      reset_n => reset_n,
      rx_clk_to_the_tse_mac => rx_clk_to_the_tse_mac,
      rx_in_to_the_fft_pipeline_0 => rx_in_to_the_fft_pipeline_0,
      set_1000_to_the_tse_mac => set_1000_to_the_tse_mac,
      set_10_to_the_tse_mac => set_10_to_the_tse_mac,
      tx_clk_to_the_tse_mac => tx_clk_to_the_tse_mac
    );


  --the_tse_mac_loopback, which is an e_instance
  the_tse_mac_loopback : tse_mac_loopback
    port map(
      gm_rx_d => gm_rx_d_to_the_tse_mac,
      gm_rx_dv => gm_rx_dv_to_the_tse_mac,
      gm_rx_err => gm_rx_err_to_the_tse_mac,
      m_rx_col => m_rx_col_to_the_tse_mac,
      m_rx_crs => m_rx_crs_to_the_tse_mac,
      m_rx_d => m_rx_d_to_the_tse_mac,
      m_rx_en => m_rx_en_to_the_tse_mac,
      m_rx_err => m_rx_err_to_the_tse_mac,
      rx_clk => rx_clk_to_the_tse_mac,
      set_10 => set_10_to_the_tse_mac,
      set_1000 => set_1000_to_the_tse_mac,
      tx_clk => tx_clk_to_the_tse_mac,
      gm_tx_d => gm_tx_d_from_the_tse_mac,
      gm_tx_en => gm_tx_en_from_the_tse_mac,
      gm_tx_err => gm_tx_err_from_the_tse_mac,
      m_tx_d => m_tx_d_from_the_tse_mac,
      m_tx_en => m_tx_en_from_the_tse_mac,
      m_tx_err => m_tx_err_from_the_tse_mac
    );


  process
  begin
    clk100MHz <= '0';
    loop
       wait for 5 ns;
       clk100MHz <= not clk100MHz;
    end loop;
  end process;
  process
  begin
    clk50Mhz <= '0';
    loop
       wait for 10 ns;
       clk50Mhz <= not clk50Mhz;
    end loop;
  end process;
  PROCESS
    BEGIN
       reset_n <= '0';
       wait for 200 ns;
       reset_n <= '1'; 
    WAIT;
  END PROCESS;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add additional architecture here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


end europa;



--synthesis translate_on
